
module dualmem(clka, clkb, dina, dinb, addra, addrb, wea, web, douta, doutb, ena, enb);

   input wire clka, clkb;
   input [7:0] dina;
   input [63:0] dinb;
   input [13:0] addra;
   input [10:0] addrb;
   input [0:0]        wea;
   input [7:0]        web;
   input [0:0]        ena, enb;
   output [7:0]       douta;
   output [63:0]      doutb;

   genvar r;

   generate for (r = 0; r < 8; r=r+1)
     RAMB16_S1_S9
     RAMB16_S1_S9_inst
       (
        .CLKA   ( clka                     ),     // Port A Clock
        .DOA    ( douta[r +: 1]            ),     // Port A 1-bit Data Output
        .ADDRA  ( addra                    ),     // Port A 14-bit Address Input
        .DIA    ( dina[r +:1]              ),     // Port A 1-bit Data Input
        .ENA    ( ena                      ),     // Port A RAM Enable Input
        .SSRA   ( 1'b0                     ),     // Port A Synchronous Set/Reset Input
        .WEA    ( wea                      ),     // Port A Write Enable Input
        .CLKB   ( clkb                     ),     // Port B Clock
        .DOB    ( doutb[r*8 +: 8]          ),     // Port B 1-bit Data Output
        .DOPB   (                          ),
        .ADDRB  ( addrb                    ),     // Port B 14-bit Address Input
        .DIB    ( dinb[r*8 +: 8]           ),     // Port B 1-bit Data Input
        .DIPB   ( 1'b0                     ),
        .ENB    ( enb                      ),     // Port B RAM Enable Input
        .SSRB   ( 1'b0                     ),     // Port B Synchronous Set/Reset Input
        .WEB    ( web[r]                   )      // Port B Write Enable Input
        );
   endgenerate

endmodule // dualmem
