// COPYRIGHT HEADER


`ifndef __UVMT_CV32_DUT_CHK_SV__
`define __UVMT_CV32_DUT_CHK_SV__


/**
 * Module encapsulating assertions for CV32 RTL DUT wrapper.
 * All ports are SV interfaces.
 */
module uvmt_cv32_dut_chk(
   uvma_debug_if  debug_if
);
   
   `pragma protect begin
   
   // TODO Add assertions to uvmt_cv32_dut_chk
   
   `pragma protect end
   
endmodule : uvmt_cv32_dut_chk


`endif // __UVMT_CV32_DUT_CHK_SV__
