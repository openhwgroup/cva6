module wt_cache_priv_adapter
  import ariane_pkg::*;
  import wt_cache_pkg::*;
  #(parameter config_pkg::cva6_cfg_t CVA6Cfg = config_pkg::cva6_cfg_empty,
    parameter type icache_areq_t = logic,
    parameter type icache_arsp_t = logic,
    parameter type icache_dreq_t = logic,
    parameter type icache_drsp_t = logic,
    parameter type dcache_req_i_t = logic,
    parameter type dcache_req_o_t = logic,
    parameter type icache_req_t = logic,
    parameter type icache_rtrn_t = logic,
    parameter int unsigned NumPorts = 4,
    parameter type noc_req_t = logic,
    parameter type noc_resp_t = logic)
   (
    input logic clk_i,
    input logic rst_ni,
    input riscv::priv_lvl_t priv_lvl_i,
    // original ports
    input logic icache_en_i,
    input logic icache_flush_i,
    output logic icache_miss_o,
    input icache_areq_t icache_areq_i,
    output icache_arsp_t icache_areq_o,
    input icache_dreq_t icache_dreq_i,
    output icache_drsp_t icache_dreq_o,
    input logic dcache_enable_i,
    input logic dcache_flush_i,
    output logic dcache_flush_ack_o,
    output logic dcache_miss_o,
    output logic [NumPorts-1:0][CVA6Cfg.DCACHE_SET_ASSOC-1:0] miss_vld_bits_o,
    input amo_req_t dcache_amo_req_i,
    output amo_resp_t dcache_amo_resp_o,
    input dcache_req_i_t [NumPorts-1:0] dcache_req_ports_i,
    output dcache_req_o_t [NumPorts-1:0] dcache_req_ports_o,
    output logic wbuffer_empty_o,
    output logic wbuffer_not_ni_o,
    output noc_req_t noc_req_o,
    input noc_resp_t noc_resp_i,
    input logic [63:0] inval_addr_i,
    input logic inval_valid_i,
    output logic inval_ready_o
   );
   // simply instantiate original subsystem, ignore priv_lvl_i
   wt_cache_subsystem #(
     .CVA6Cfg(CVA6Cfg),
     .icache_areq_t(icache_areq_t),
     .icache_arsp_t(icache_arsp_t),
     .icache_dreq_t(icache_dreq_t),
     .icache_drsp_t(icache_drsp_t),
     .dcache_req_i_t(dcache_req_i_t),
     .dcache_req_o_t(dcache_req_o_t),
     .icache_req_t(icache_req_t),
     .icache_rtrn_t(icache_rtrn_t),
     .NumPorts(NumPorts),
     .noc_req_t(noc_req_t),
     .noc_resp_t(noc_resp_t)
   ) i_wt_cache_subsystem (
     .clk_i(clk_i),
     .rst_ni(rst_ni),
     .icache_en_i(icache_en_i),
     .icache_flush_i(icache_flush_i),
     .icache_miss_o(icache_miss_o),
     .icache_areq_i(icache_areq_i),
     .icache_areq_o(icache_areq_o),
     .icache_dreq_i(icache_dreq_i),
     .icache_dreq_o(icache_dreq_o),
     .dcache_enable_i(dcache_enable_i),
     .dcache_flush_i(dcache_flush_i),
     .dcache_flush_ack_o(dcache_flush_ack_o),
     .dcache_miss_o(dcache_miss_o),
     .miss_vld_bits_o(miss_vld_bits_o),
     .dcache_amo_req_i(dcache_amo_req_i),
     .dcache_amo_resp_o(dcache_amo_resp_o),
     .dcache_req_ports_i(dcache_req_ports_i),
     .dcache_req_ports_o(dcache_req_ports_o),
     .wbuffer_empty_o(wbuffer_empty_o),
     .wbuffer_not_ni_o(wbuffer_not_ni_o),
     .noc_req_o(noc_req_o),
     .noc_resp_i(noc_resp_i),
     .inval_addr_i(inval_addr_i),
     .inval_valid_i(inval_valid_i),
     .inval_ready_o(inval_ready_o)
   );
endmodule
