// Copyright 2020 OpenHW Group
// Copyright 2020 Datum Technology Corporation
// Copyright 2020 Silicon Labs, Inc.
//
// Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// 
//     https://solderpad.org/licenses/
// 
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


`ifndef __UVMA_ISACOV_MACROS_SV__
`define __UVMA_ISACOV_MACROS_SV__


`define ISACOV_CP_BITWISE(name, field, iff_exp) \
``name``: coverpoint(``field``) iff (``iff_exp``) { \
    wildcard bins BIT0_0  = {32'b???????????????????????????????0}; \
    wildcard bins BIT1_0  = {32'b??????????????????????????????0?}; \
    wildcard bins BIT2_0  = {32'b?????????????????????????????0??}; \
    wildcard bins BIT3_0  = {32'b????????????????????????????0???}; \
    wildcard bins BIT4_0  = {32'b???????????????????????????0????}; \
    wildcard bins BIT5_0  = {32'b??????????????????????????0?????}; \
    wildcard bins BIT6_0  = {32'b?????????????????????????0??????}; \
    wildcard bins BIT7_0  = {32'b????????????????????????0???????}; \
    wildcard bins BIT8_0  = {32'b???????????????????????0????????}; \
    wildcard bins BIT9_0  = {32'b??????????????????????0?????????}; \
    wildcard bins BIT10_0 = {32'b?????????????????????0??????????}; \
    wildcard bins BIT11_0 = {32'b????????????????????0???????????}; \
    wildcard bins BIT12_0 = {32'b???????????????????0????????????}; \
    wildcard bins BIT13_0 = {32'b??????????????????0?????????????}; \
    wildcard bins BIT14_0 = {32'b?????????????????0??????????????}; \
    wildcard bins BIT15_0 = {32'b????????????????0???????????????}; \
    wildcard bins BIT16_0 = {32'b???????????????0????????????????}; \
    wildcard bins BIT17_0 = {32'b??????????????0?????????????????}; \
    wildcard bins BIT18_0 = {32'b?????????????0??????????????????}; \
    wildcard bins BIT19_0 = {32'b????????????0???????????????????}; \
    wildcard bins BIT20_0 = {32'b???????????0????????????????????}; \
    wildcard bins BIT21_0 = {32'b??????????0?????????????????????}; \
    wildcard bins BIT22_0 = {32'b?????????0??????????????????????}; \
    wildcard bins BIT23_0 = {32'b????????0???????????????????????}; \
    wildcard bins BIT24_0 = {32'b???????0????????????????????????}; \
    wildcard bins BIT25_0 = {32'b??????0?????????????????????????}; \
    wildcard bins BIT26_0 = {32'b?????0??????????????????????????}; \
    wildcard bins BIT27_0 = {32'b????0???????????????????????????}; \
    wildcard bins BIT28_0 = {32'b???0????????????????????????????}; \
    wildcard bins BIT29_0 = {32'b??0?????????????????????????????}; \
    wildcard bins BIT30_0 = {32'b?0??????????????????????????????}; \
    wildcard bins BIT31_0 = {32'b0???????????????????????????????}; \
    wildcard bins BIT0_1  = {32'b???????????????????????????????1}; \
    wildcard bins BIT1_1  = {32'b??????????????????????????????1?}; \
    wildcard bins BIT2_1  = {32'b?????????????????????????????1??}; \
    wildcard bins BIT3_1  = {32'b????????????????????????????1???}; \
    wildcard bins BIT4_1  = {32'b???????????????????????????1????}; \
    wildcard bins BIT5_1  = {32'b??????????????????????????1?????}; \
    wildcard bins BIT6_1  = {32'b?????????????????????????1??????}; \
    wildcard bins BIT7_1  = {32'b????????????????????????1???????}; \
    wildcard bins BIT8_1  = {32'b???????????????????????1????????}; \
    wildcard bins BIT9_1  = {32'b??????????????????????1?????????}; \
    wildcard bins BIT10_1 = {32'b?????????????????????1??????????}; \
    wildcard bins BIT11_1 = {32'b????????????????????1???????????}; \
    wildcard bins BIT12_1 = {32'b???????????????????1????????????}; \
    wildcard bins BIT13_1 = {32'b??????????????????1?????????????}; \
    wildcard bins BIT14_1 = {32'b?????????????????1??????????????}; \
    wildcard bins BIT15_1 = {32'b????????????????1???????????????}; \
    wildcard bins BIT16_1 = {32'b???????????????1????????????????}; \
    wildcard bins BIT17_1 = {32'b??????????????1?????????????????}; \
    wildcard bins BIT18_1 = {32'b?????????????1??????????????????}; \
    wildcard bins BIT19_1 = {32'b????????????1???????????????????}; \
    wildcard bins BIT20_1 = {32'b???????????1????????????????????}; \
    wildcard bins BIT21_1 = {32'b??????????1?????????????????????}; \
    wildcard bins BIT22_1 = {32'b?????????1??????????????????????}; \
    wildcard bins BIT23_1 = {32'b????????1???????????????????????}; \
    wildcard bins BIT24_1 = {32'b???????1????????????????????????}; \
    wildcard bins BIT25_1 = {32'b??????1?????????????????????????}; \
    wildcard bins BIT26_1 = {32'b?????1??????????????????????????}; \
    wildcard bins BIT27_1 = {32'b????1???????????????????????????}; \
    wildcard bins BIT28_1 = {32'b???1????????????????????????????}; \
    wildcard bins BIT29_1 = {32'b??1?????????????????????????????}; \
    wildcard bins BIT30_1 = {32'b?1??????????????????????????????}; \
    wildcard bins BIT31_1 = {32'b1???????????????????????????????}; \
}

`define ISACOV_CP_BITWISE_31_12(name, field, iff_exp) \
``name``: coverpoint(``field``) iff (``iff_exp``) { \
    wildcard bins BIT12_0 = {32'b???????????????????0????????????}; \
    wildcard bins BIT13_0 = {32'b??????????????????0?????????????}; \
    wildcard bins BIT14_0 = {32'b?????????????????0??????????????}; \
    wildcard bins BIT15_0 = {32'b????????????????0???????????????}; \
    wildcard bins BIT16_0 = {32'b???????????????0????????????????}; \
    wildcard bins BIT17_0 = {32'b??????????????0?????????????????}; \
    wildcard bins BIT18_0 = {32'b?????????????0??????????????????}; \
    wildcard bins BIT19_0 = {32'b????????????0???????????????????}; \
    wildcard bins BIT20_0 = {32'b???????????0????????????????????}; \
    wildcard bins BIT21_0 = {32'b??????????0?????????????????????}; \
    wildcard bins BIT22_0 = {32'b?????????0??????????????????????}; \
    wildcard bins BIT23_0 = {32'b????????0???????????????????????}; \
    wildcard bins BIT24_0 = {32'b???????0????????????????????????}; \
    wildcard bins BIT25_0 = {32'b??????0?????????????????????????}; \
    wildcard bins BIT26_0 = {32'b?????0??????????????????????????}; \
    wildcard bins BIT27_0 = {32'b????0???????????????????????????}; \
    wildcard bins BIT28_0 = {32'b???0????????????????????????????}; \
    wildcard bins BIT29_0 = {32'b??0?????????????????????????????}; \
    wildcard bins BIT30_0 = {32'b?0??????????????????????????????}; \
    wildcard bins BIT31_0 = {32'b0???????????????????????????????}; \
    wildcard bins BIT12_1 = {32'b???????????????????1????????????}; \
    wildcard bins BIT13_1 = {32'b??????????????????1?????????????}; \
    wildcard bins BIT14_1 = {32'b?????????????????1??????????????}; \
    wildcard bins BIT15_1 = {32'b????????????????1???????????????}; \
    wildcard bins BIT16_1 = {32'b???????????????1????????????????}; \
    wildcard bins BIT17_1 = {32'b??????????????1?????????????????}; \
    wildcard bins BIT18_1 = {32'b?????????????1??????????????????}; \
    wildcard bins BIT19_1 = {32'b????????????1???????????????????}; \
    wildcard bins BIT20_1 = {32'b???????????1????????????????????}; \
    wildcard bins BIT21_1 = {32'b??????????1?????????????????????}; \
    wildcard bins BIT22_1 = {32'b?????????1??????????????????????}; \
    wildcard bins BIT23_1 = {32'b????????1???????????????????????}; \
    wildcard bins BIT24_1 = {32'b???????1????????????????????????}; \
    wildcard bins BIT25_1 = {32'b??????1?????????????????????????}; \
    wildcard bins BIT26_1 = {32'b?????1??????????????????????????}; \
    wildcard bins BIT27_1 = {32'b????1???????????????????????????}; \
    wildcard bins BIT28_1 = {32'b???1????????????????????????????}; \
    wildcard bins BIT29_1 = {32'b??1?????????????????????????????}; \
    wildcard bins BIT30_1 = {32'b?1??????????????????????????????}; \
    wildcard bins BIT31_1 = {32'b1???????????????????????????????}; \
} \

`define ISACOV_CP_BITWISE_19_0(name, field, iff_exp) \
``name``: coverpoint(``field``) iff (``iff_exp``) { \
    wildcard bins BIT0_0  = {20'b???????????????????0}; \
    wildcard bins BIT1_0  = {20'b??????????????????0?}; \
    wildcard bins BIT2_0  = {20'b?????????????????0??}; \
    wildcard bins BIT3_0  = {20'b????????????????0???}; \
    wildcard bins BIT4_0  = {20'b???????????????0????}; \
    wildcard bins BIT5_0  = {20'b??????????????0?????}; \
    wildcard bins BIT6_0  = {20'b?????????????0??????}; \
    wildcard bins BIT7_0  = {20'b????????????0???????}; \
    wildcard bins BIT8_0  = {20'b???????????0????????}; \
    wildcard bins BIT9_0  = {20'b??????????0?????????}; \
    wildcard bins BIT10_0 = {20'b?????????0??????????}; \
    wildcard bins BIT11_0 = {20'b????????0???????????}; \
    wildcard bins BIT12_0 = {20'b???????0????????????}; \
    wildcard bins BIT13_0 = {20'b??????0?????????????}; \
    wildcard bins BIT14_0 = {20'b?????0??????????????}; \
    wildcard bins BIT15_0 = {20'b????0???????????????}; \
    wildcard bins BIT16_0 = {20'b???0????????????????}; \
    wildcard bins BIT17_0 = {20'b??0?????????????????}; \
    wildcard bins BIT18_0 = {20'b?0??????????????????}; \
    wildcard bins BIT19_0 = {20'b0???????????????????}; \
    wildcard bins BIT0_1  = {20'b???????????????????1}; \
    wildcard bins BIT1_1  = {20'b??????????????????1?}; \
    wildcard bins BIT2_1  = {20'b?????????????????1??}; \
    wildcard bins BIT3_1  = {20'b????????????????1???}; \
    wildcard bins BIT4_1  = {20'b???????????????1????}; \
    wildcard bins BIT5_1  = {20'b??????????????1?????}; \
    wildcard bins BIT6_1  = {20'b?????????????1??????}; \
    wildcard bins BIT7_1  = {20'b????????????1???????}; \
    wildcard bins BIT8_1  = {20'b???????????1????????}; \
    wildcard bins BIT9_1  = {20'b??????????1?????????}; \
    wildcard bins BIT10_1 = {20'b?????????1??????????}; \
    wildcard bins BIT11_1 = {20'b????????1???????????}; \
    wildcard bins BIT12_1 = {20'b???????1????????????}; \
    wildcard bins BIT13_1 = {20'b??????1?????????????}; \
    wildcard bins BIT14_1 = {20'b?????1??????????????}; \
    wildcard bins BIT15_1 = {20'b????1???????????????}; \
    wildcard bins BIT16_1 = {20'b???1????????????????}; \
    wildcard bins BIT17_1 = {20'b??1?????????????????}; \
    wildcard bins BIT18_1 = {20'b?1??????????????????}; \
    wildcard bins BIT19_1 = {20'b1???????????????????}; \
}

`define ISACOV_CP_BITWISE_11_0(name, field, iff_exp) \
``name``: coverpoint(``field``) iff (``iff_exp``) { \
    wildcard bins BIT0_0  = {12'b???????????0}; \
    wildcard bins BIT1_0  = {12'b??????????0?}; \
    wildcard bins BIT2_0  = {12'b?????????0??}; \
    wildcard bins BIT3_0  = {12'b????????0???}; \
    wildcard bins BIT4_0  = {12'b???????0????}; \
    wildcard bins BIT5_0  = {12'b??????0?????}; \
    wildcard bins BIT6_0  = {12'b?????0??????}; \
    wildcard bins BIT7_0  = {12'b????0???????}; \
    wildcard bins BIT8_0  = {12'b???0????????}; \
    wildcard bins BIT9_0  = {12'b??0?????????}; \
    wildcard bins BIT10_0 = {12'b?0??????????}; \
    wildcard bins BIT11_0 = {12'b0???????????}; \
    wildcard bins BIT0_1  = {12'b???????????1}; \
    wildcard bins BIT1_1  = {12'b??????????1?}; \
    wildcard bins BIT2_1  = {12'b?????????1??}; \
    wildcard bins BIT3_1  = {12'b????????1???}; \
    wildcard bins BIT4_1  = {12'b???????1????}; \
    wildcard bins BIT5_1  = {12'b??????1?????}; \
    wildcard bins BIT6_1  = {12'b?????1??????}; \
    wildcard bins BIT7_1  = {12'b????1???????}; \
    wildcard bins BIT8_1  = {12'b???1????????}; \
    wildcard bins BIT9_1  = {12'b??1?????????}; \
    wildcard bins BIT10_1 = {12'b?1??????????}; \
    wildcard bins BIT11_1 = {12'b1???????????}; \
}

`endif // __UVMA_ISACOV_MACROS_SV__
