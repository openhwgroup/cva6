`define NEXYS_VIDEO

`define ARIANE_DATA_WIDTH 64

// Instantiate protocol checker
// `define PROTOCOL_CHECKER

// write-back cache
// `define WB_DCACHE

// write-through cache
`define WT_DCACHE

`define RAMB16
