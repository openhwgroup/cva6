riscv_CV32E40P.sv