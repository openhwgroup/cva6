// COPYRIGHT HEADER


`ifndef __UVMA_DEBUG_MACROS_SV__
`define __UVMA_DEBUG_MACROS_SV__





`endif // __UVMA_DEBUG_MACROS_SV__
