// COPYRIGHT HEADER


`ifndef __UVML_TRN_TDEFS_SV__
`define __UVML_TRN_TDEFS_SV__





`endif // __UVML_TRN_TDEFS_SV__
