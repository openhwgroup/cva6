// COPYRIGHT HEADER


`ifndef __UVMT_CV32_TDEFS_SV__
`define __UVMT_CV32_TDEFS_SV__





`endif // __UVMT_CV32_TDEFS_SV__
