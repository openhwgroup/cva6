/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the “License”); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 216;

    const logic [RomSize-1:0][63:0] mem = {
        64'h006b_636f6c63,
        64'h00737470_75727265,
        64'h746e6900_746e6572,
        64'h61702d74_70757272,
        64'h65746e69_00766564,
        64'h6e2c7663_73697200,
        64'h79746972_6f697270,
        64'h2d78616d_2c766373,
        64'h69720073_656d616e,
        64'h2d676572_00646564,
        64'h6e657478_652d7374,
        64'h70757272_65746e69,
        64'h00736567_6e617200,
        64'h656c646e_6168702c,
        64'h78756e69_6c007265,
        64'h6c6c6f72_746e6f63,
        64'h2d747075_72726574,
        64'h6e690073_6c6c6563,
        64'h2d747075_72726574,
        64'h6e692300_79636e65,
        64'h75716572_662d6b63,
        64'h6f6c6300_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h006c6564_6f6d0065,
        64'h6c626974_61706d6f,
        64'h6300736c_6c65632d,
        64'h657a6973_2300736c,
        64'h6c65632d_73736572,
        64'h64646123_09000000,
        64'h02000000_02000000,
        64'h00000030_66697468,
        64'h2c626375_1b000000,
        64'h0a000000_03000000,
        64'h00000000_66697468,
        64'h01000000_02000000,
        64'h02000000_80f0fa02,
        64'h0c010000_04000000,
        64'h03000000_02000000,
        64'h01000000_00000000,
        64'h01010000_0c000000,
        64'h03000000_02000000,
        64'hf0000000_04000000,
        64'h03000000_00000100,
        64'h00000000_00000010,
        64'h00000000_4b000000,
        64'h10000000_03000000,
        64'h00000000_612e3230,
        64'h2e312d65_74696c74,
        64'h7261752d_6978612c,
        64'h786e6c78_1b000000,
        64'h19000000_03000000,
        64'h00000030_30303030,
        64'h30303140_74726175,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'hc8000000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000000,
        64'h00000000_4b000000,
        64'h10000000_03000000,
        64'hffff0000_01000000,
        64'hb4000000_08000000,
        64'h03000000_00333130,
        64'h2d677562_65642c76,
        64'h63736972_1b000000,
        64'h10000000_03000000,
        64'h00003040_72656c6c,
        64'h6f72746e_6f632d67,
        64'h75626564_01000000,
        64'h02000000_02000000,
        64'ha5000000_04000000,
        64'h03000000_02000000,
        64'h9f000000_04000000,
        64'h03000000_02000000,
        64'he5000000_04000000,
        64'h03000000_07000000,
        64'hd2000000_04000000,
        64'h03000000_006c6f72,
        64'h746e6f63_c8000000,
        64'h08000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h4b000000_10000000,
        64'h03000000_09000000,
        64'h01000000_0b000000,
        64'h01000000_b4000000,
        64'h10000000_03000000,
        64'h8a000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h79000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_00000c00,
        64'h00000000_00000002,
        64'h00000000_4b000000,
        64'h10000000_03000000,
        64'h07000000_01000000,
        64'h03000000_01000000,
        64'hb4000000_10000000,
        64'h03000000_00000000,
        64'h30746e69_6c632c76,
        64'h63736972_1b000000,
        64'h0d000000_03000000,
        64'h00000030_30303030,
        64'h30324074_6e696c63,
        64'h01000000_ad000000,
        64'h00000000_03000000,
        64'h00007375_622d656c,
        64'h706d6973_00636f73,
        64'h2d657261_622d656e,
        64'h61697261_2c687465,
        64'h1b000000_1f000000,
        64'h03000000_02000000,
        64'h0f000000_04000000,
        64'h03000000_02000000,
        64'h00000000_04000000,
        64'h03000000_00636f73,
        64'h01000000_02000000,
        64'h00000002_00000000,
        64'h00000080_00000000,
        64'h4b000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_3f000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h01000000_a5000000,
        64'h04000000_03000000,
        64'h01000000_9f000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_8a000000,
        64'h00000000_03000000,
        64'h01000000_79000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_80f0fa02,
        64'h69000000_04000000,
        64'h03000000_00003933,
        64'h76732c76_63736972,
        64'h60000000_0b000000,
        64'h03000000_00000000,
        64'h63616d69_34367672,
        64'h56000000_09000000,
        64'h03000000_00000076,
        64'h63736972_1b000000,
        64'h06000000_03000000,
        64'h00000000_79616b6f,
        64'h4f000000_05000000,
        64'h03000000_00000000,
        64'h4b000000_04000000,
        64'h03000000_00757063,
        64'h3f000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_2c000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hf4040000_12010000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h2c050000_38000000,
        64'h3e060000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_0000bff5,
        64'h10500073_03c58593,
        64'h00000597_f1402573,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00008402_07458593,
        64'h00000597_f1402573,
        64'h01f41413_0010041b
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    assign rdata_o = mem[addr_q];
endmodule
