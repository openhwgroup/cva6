// COPYRIGHT HEADER


`ifndef __UVML_HRTBT_MACROS_SV__
`define __UVML_HRTBT_MACROS_SV__


`define uvml_hrtbt(ID)
`define uvml_hrtbt_set_cfg(NAME, VALUE)


`endif // __UVML_HRTBT_MACROS_SV__
