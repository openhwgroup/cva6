// COPYRIGHT HEADER


`ifndef __UVMA_DEBUG_IF_CHK_SV__
`define __UVMA_DEBUG_IF_CHK_SV__


/**
 * Encapsulates assertions targeting uvma_debug_if.
 */
module uvma_debug_if_chk(
   uvma_debug_if  debug_if
);
   
   `pragma protect begin
   
   // TODO Add assertions to uvma_debug_if_chk
   
   `pragma protect end
   
endmodule : uvma_debug_if_chk


`endif // __UVMA_DEBUG_IF_CHK_SV__
