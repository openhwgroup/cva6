// Copyright 2021 Thales DIS design services SAS
//
// Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.0
// You may obtain a copy of the License at https://solderpad.org/licenses/
//
// Original Author: Zineb EL KACIMI (zineb.el-kacimi@external.thalesgroup.com)


`ifndef __UVMA_CVXIF_CONSTANTS_SV__
`define __UVMA_CVXIF_CONSTANTS_SV__


const int unsigned  uvma_cvxif_issue_ready_min     = 4;
const int unsigned  uvma_cvxif_issue_ready_max     = 10;
const int unsigned  uvma_cvxif_issue_not_ready_min = 1;
const int unsigned  uvma_cvxif_issue_not_ready_max = 2;


`endif //__UVMA_CVXIF_CONSTANTS_SV__
