class reset_sequence extends fu_if_seq;

   `uvm_object_utils(reset_sequence);

   function new(string name = "reset");
      super.new(name);
   endfunction : new


   task body();
      
      fu_if_seq_item command;

      command = fu_if_seq_item::type_id::create("command");
      `uvm_info("RESET", "Starting reset phase", UVM_MEDIUM);
      // reset 
      for (int i = 0; i < 20; i++) begin
      start_item(command);
      command.operand_a = 0;
      command.operand_b = 0;
      command.operand_c = 0;
      command.operator = 7'b00;
      finish_item(command);
      end

   endtask : body
endclass : reset_sequence
