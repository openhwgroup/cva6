// COPYRIGHT HEADER


`ifndef __UVMA_RESET_CONSTANTS_SV__
`define __UVMA_RESET_CONSTANTS_SV__





`endif // __UVMA_RESET_CONSTANTS_SV__
