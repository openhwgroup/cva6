// Copyright 2018 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

// Xilinx FPGA top-level
module ariane_xilinx (
`ifdef VCU118
  input  wire          c0_sys_clk_p    ,  // 250 MHz Clock for DDR
  input  wire          c0_sys_clk_n    ,  // 250 MHz Clock for DDR
  input  wire          sys_clk_p       ,  // 100 MHz Clock for PCIe
  input  wire          sys_clk_n       ,  // 100 MHz Clock for PCIE
  input  wire          sys_rst_n       ,  // PCIe Reset
  input  logic         cpu_reset       ,  // CPU subsystem reset
  output wire [16 : 0] c0_ddr4_adr     ,
  output wire [1 : 0]  c0_ddr4_ba      ,
  output wire [0 : 0]  c0_ddr4_cke     ,
  output wire [0 : 0]  c0_ddr4_cs_n    ,
  inout  wire [7 : 0]  c0_ddr4_dm_dbi_n,
  inout  wire [63 : 0] c0_ddr4_dq      ,
  inout  wire [7 : 0]  c0_ddr4_dqs_c   ,
  inout  wire [7 : 0]  c0_ddr4_dqs_t   ,
  output wire [0 : 0]  c0_ddr4_odt     ,
  output wire [0 : 0]  c0_ddr4_bg      ,
  output wire          c0_ddr4_reset_n ,
  output wire          c0_ddr4_act_n   ,
  output wire [0 : 0]  c0_ddr4_ck_c    ,
  output wire [0 : 0]  c0_ddr4_ck_t    ,
  output wire [7 : 0]  pci_exp_txp     ,
  output wire [7 : 0]  pci_exp_txn     ,
  input  wire [7 : 0]  pci_exp_rxp     ,
  input  wire [7 : 0]  pci_exp_rxn     ,
`elsif GENESYSII
  input  logic         sys_clk_p   ,
  input  logic         sys_clk_n   ,
  input  logic         cpu_resetn  ,
  inout  logic [31:0]  ddr3_dq     ,
  inout  logic [ 3:0]  ddr3_dqs_n  ,
  inout  logic [ 3:0]  ddr3_dqs_p  ,
  output logic [14:0]  ddr3_addr   ,
  output logic [ 2:0]  ddr3_ba     ,
  output logic         ddr3_ras_n  ,
  output logic         ddr3_cas_n  ,
  output logic         ddr3_we_n   ,
  output logic         ddr3_reset_n,
  output logic [ 0:0]  ddr3_ck_p   ,
  output logic [ 0:0]  ddr3_ck_n   ,
  output logic [ 0:0]  ddr3_cke    ,
  output logic [ 0:0]  ddr3_cs_n   ,
  output logic [ 3:0]  ddr3_dm     ,
  output logic [ 0:0]  ddr3_odt    ,
  output logic [ 7:0]  led         ,
  input  logic [ 7:0]  sw          ,
  output logic         fan_pwm     ,
`endif
  // SPI
  output logic        spi_mosi    ,
  input  logic        spi_miso    ,
  output logic        spi_ss      ,
  output logic        spi_clk_o   ,
  output logic        spi_mosi_2  ,
  output logic        spi_miso_2  ,
  output logic        spi_ss_2    ,
  output logic        spi_clk_o_2 ,
  // common part
  input  logic        tck         ,
  input  logic        tms         ,
  input  logic        trst_n      ,
  input  logic        tdi         ,
  output logic        tdo         ,
  input  logic        rx          ,
  output logic        tx
);
// 24 MByte in 8 byte words
localparam NumWords = (24 * 1024 * 1024) / 8;
localparam NBSlave = 4; // debug, Instruction fetch, data bypass, data
localparam CacheStartAddr = (1 << 31);
localparam AxiAddrWidth = 64;
localparam AxiDataWidth = 64;
localparam AxiIdWidthMaster = 2;
localparam AxiIdWidthSlaves = AxiIdWidthMaster + $clog2(NBSlave); // 4
localparam AxiUserWidth = 1;

AXI_BUS #(
    .AXI_ADDR_WIDTH ( AxiAddrWidth     ),
    .AXI_DATA_WIDTH ( AxiDataWidth     ),
    .AXI_ID_WIDTH   ( AxiIdWidthMaster ),
    .AXI_USER_WIDTH ( AxiUserWidth     )
) slave[NBSlave-1:0]();

AXI_BUS #(
    .AXI_ADDR_WIDTH ( AxiAddrWidth     ),
    .AXI_DATA_WIDTH ( AxiDataWidth     ),
    .AXI_ID_WIDTH   ( AxiIdWidthMaster ),
    .AXI_USER_WIDTH ( AxiUserWidth     )
) dummy_slave();

AXI_BUS #(
    .AXI_ADDR_WIDTH ( AxiAddrWidth     ),
    .AXI_DATA_WIDTH ( AxiDataWidth     ),
    .AXI_ID_WIDTH   ( AxiIdWidthMaster ),
    .AXI_USER_WIDTH ( AxiUserWidth     )
) slave_slice[NBSlave-1:0]();

AXI_BUS #(
    .AXI_ADDR_WIDTH ( AxiAddrWidth     ),
    .AXI_DATA_WIDTH ( AxiDataWidth     ),
    .AXI_ID_WIDTH   ( AxiIdWidthSlaves ),
    .AXI_USER_WIDTH ( AxiUserWidth     )
) master[ariane_soc::NB_PERIPHERALS-1:0]();

// spi hack
assign spi_mosi_2 = spi_mosi;
assign spi_miso_2 = spi_miso;
assign spi_clk_o_2 = spi_clk_o;
assign spi_ss_2 = spi_ss;

// disable test-enable
logic test_en;
logic ndmreset;
logic ndmreset_n;
logic debug_req_irq;
logic time_irq;
logic ipi;

logic clk;
logic spi_clk_i;
logic ddr_sync_reset;
logic ddr_clock_out;

logic rst_n, rst;
logic rtc;

// we need to switch reset polarity
`ifdef VCU118
logic cpu_resetn;
assign cpu_resetn = ~cpu_reset;
`elsif GENESYSII
logic cpu_reset;
assign cpu_reset  = ~cpu_resetn;
`endif

assign rst_n      = ~ddr_sync_reset;
assign rst        = ddr_sync_reset;

// ROM
logic                    rom_req;
logic [AxiAddrWidth-1:0] rom_addr;
logic [AxiDataWidth-1:0] rom_rdata;

// Debug
logic          debug_req_valid;
logic          debug_req_ready;
dm::dmi_req_t  debug_req;
logic          debug_resp_valid;
logic          debug_resp_ready;
dm::dmi_resp_t debug_resp;

logic dmactive;

// IRQ
logic [1:0] irq;
assign test_en    = 1'b0;
assign ndmreset_n = ~ndmreset ;

logic [NBSlave-1:0] pc_asserted;

// Slice the AXI Masters (slave ports on the XBar)
for (genvar i = 0; i < NBSlave; i++) begin : slave_cut_gen
    axi_cut #(
        .ADDR_WIDTH ( AxiAddrWidth     ),
        .DATA_WIDTH ( AxiDataWidth     ),
        .ID_WIDTH   ( AxiIdWidthMaster ),
        .USER_WIDTH ( AxiUserWidth     )
    ) i_axi_cut (
        .clk_i  ( clk            ),
        .rst_ni ( ndmreset_n     ),
        .in     ( slave_slice[i] ),
        .out    ( slave[i]       )
    );

    if (ariane_soc::GenProtocolChecker) begin : gen_protocol_check
      axi_protocol_checker_0 i_axi_protocol_checker (
        .pc_status( ), // debug probe
        .pc_asserted(pc_asserted[i]),
        .aclk(clk),
        .aresetn(ndmreset_n),
        .pc_axi_awid(slave[i].aw_id),
        .pc_axi_awaddr(slave[i].aw_addr),
        .pc_axi_awlen(slave[i].aw_len),
        .pc_axi_awsize(slave[i].aw_size),
        .pc_axi_awburst(slave[i].aw_burst),
        .pc_axi_awlock(slave[i].aw_lock),
        .pc_axi_awcache(slave[i].aw_cache),
        .pc_axi_awprot(slave[i].aw_prot),
        .pc_axi_awqos(slave[i].aw_qos),
        .pc_axi_awregion(slave[i].aw_region),
        .pc_axi_awready(slave[i].aw_ready),
        .pc_axi_awvalid(slave[i].aw_valid),
        .pc_axi_awuser(slave[i].aw_user),
        .pc_axi_wlast(slave[i].w_last),
        .pc_axi_wdata(slave[i].w_data),
        .pc_axi_wstrb(slave[i].w_strb),
        .pc_axi_wuser(slave[i].w_user),
        .pc_axi_wvalid(slave[i].w_valid),
        .pc_axi_wready(slave[i].w_ready),
        .pc_axi_bid(slave[i].b_id),
        .pc_axi_bresp(slave[i].b_resp),
        .pc_axi_buser(slave[i].b_user),
        .pc_axi_bvalid(slave[i].b_valid),
        .pc_axi_bready(slave[i].b_ready),
        .pc_axi_arid(slave[i].ar_id),
        .pc_axi_araddr(slave[i].ar_addr),
        .pc_axi_arlen(slave[i].ar_len),
        .pc_axi_arsize(slave[i].ar_size),
        .pc_axi_arburst(slave[i].ar_burst),
        .pc_axi_arlock(slave[i].ar_lock),
        .pc_axi_arcache(slave[i].ar_cache),
        .pc_axi_arprot(slave[i].ar_prot),
        .pc_axi_arqos(slave[i].ar_qos),
        .pc_axi_arregion(slave[i].ar_region),
        .pc_axi_aruser(slave[i].ar_user),
        .pc_axi_arvalid(slave[i].ar_valid),
        .pc_axi_arready(slave[i].ar_ready),
        .pc_axi_rid(slave[i].r_id),
        .pc_axi_rlast(slave[i].r_last),
        .pc_axi_rdata(slave[i].r_data),
        .pc_axi_rresp(slave[i].r_resp),
        .pc_axi_ruser(slave[i].r_user),
        .pc_axi_rvalid(slave[i].r_valid),
        .pc_axi_rready(slave[i].r_ready)
      );
    end
end

// ---------------
// AXI Xbar
// ---------------
axi_node_wrap_with_slices #(
    // three ports from Ariane (instruction, data and bypass)
    .NB_SLAVE           ( NBSlave                    ),
    .NB_MASTER          ( ariane_soc::NB_PERIPHERALS ),
    .AXI_ADDR_WIDTH     ( AxiAddrWidth               ),
    .AXI_DATA_WIDTH     ( AxiDataWidth               ),
    .AXI_USER_WIDTH     ( AxiUserWidth               ),
    .AXI_ID_WIDTH       ( AxiIdWidthMaster           ),
    .MASTER_SLICE_DEPTH ( 2                          ),
    .SLAVE_SLICE_DEPTH  ( 2                          )
) i_axi_xbar (
    .clk          ( clk        ),
    .rst_n        ( ndmreset_n ),
    .test_en_i    ( test_en    ),
    .slave        ( slave      ),
    .master       ( master     ),
    .start_addr_i ({
        ariane_soc::DebugBase,
        ariane_soc::ROMBase,
        ariane_soc::CLINTBase,
        ariane_soc::PLICBase,
        ariane_soc::UARTBase,
        ariane_soc::SPIBase,
`ifdef INCL_SRAM
        ariane_soc::SRAMBase,
        ariane_soc::DRAMBase
`else
        ariane_soc::DRAMBase
`endif
    }),
    .end_addr_i   ({
        ariane_soc::DebugBase + ariane_soc::DebugLength - 1,
        ariane_soc::ROMBase   + ariane_soc::ROMLength - 1,
        ariane_soc::CLINTBase + ariane_soc::CLINTLength - 1,
        ariane_soc::PLICBase  + ariane_soc::PLICLength - 1,
        ariane_soc::UARTBase  + ariane_soc::UARTLength - 1,
        ariane_soc::SPIBase   + ariane_soc::SPILength - 1,
`ifdef INCL_SRAM
        ariane_soc::SRAMBase  + ariane_soc::SRAMLength - 1,
        ariane_soc::DRAMBase  + ariane_soc::DRAMLength - 1
`else
        ariane_soc::DRAMBase  + ariane_soc::DRAMLength - 1
`endif
    })
);

// ---------------
// Debug Module
// ---------------
dmi_jtag i_dmi_jtag (
    .clk_i                ( clk                  ),
    .rst_ni               ( rst_n                ),
    .dmi_rst_no           (                      ), // keep open
    .dmi_req_valid_o      ( debug_req_valid      ),
    .dmi_req_ready_i      ( debug_req_ready      ),
    .dmi_req_o            ( debug_req            ),
    .dmi_resp_valid_i     ( debug_resp_valid     ),
    .dmi_resp_ready_o     ( debug_resp_ready     ),
    .dmi_resp_i           ( debug_resp           ),
    .tck_i                ( tck    ),
    .tms_i                ( tms    ),
    .trst_ni              ( trst_n ),
    .td_i                 ( tdi    ),
    .td_o                 ( tdo    ),
    .tdo_oe_o             (        )
);

// debug module
dm_top #(
    // current implementation only supports 1 hart
    .NrHarts              ( 1                    ),
    .AxiIdWidth           ( AxiIdWidthSlaves     ),
    .AxiAddrWidth         ( AxiAddrWidth         ),
    .AxiDataWidth         ( AxiDataWidth         ),
    .AxiUserWidth         ( AxiUserWidth         )
) i_dm_top (
    .clk_i                ( clk                        ),
    .rst_ni               ( rst_n                      ), // PoR
    .testmode_i           ( test_en                    ),
    .ndmreset_o           ( ndmreset                   ),
    .dmactive_o           ( dmactive                   ), // active debug session
    .debug_req_o          ( debug_req_irq              ),
    .unavailable_i        ( '0                         ),
    .axi_master           ( dummy_slave                ),
    .axi_slave            ( master[ariane_soc::Debug]  ),
    .dmi_rst_ni           ( rst_n                      ),
    .dmi_req_valid_i      ( debug_req_valid            ),
    .dmi_req_ready_o      ( debug_req_ready            ),
    .dmi_req_i            ( debug_req                  ),
    .dmi_resp_valid_o     ( debug_resp_valid           ),
    .dmi_resp_ready_i     ( debug_resp_ready           ),
    .dmi_resp_o           ( debug_resp                 )
);

assign dummy_slave.aw_ready = 1'b0;
assign dummy_slave.ar_ready = 1'b0;
assign dummy_slave.w_ready = 1'b0;
assign dummy_slave.b_valid = 1'b0;
assign dummy_slave.r_valid = 1'b0;

// ---------------
// Core
// ---------------
ariane #(
    .CACHE_START_ADDR ( CacheStartAddr   ),
    .AXI_ID_WIDTH     ( AxiIdWidthMaster ),
    .AXI_USER_WIDTH   ( AxiUserWidth     )
) i_ariane (
    .clk_i                ( clk                 ),
    .rst_ni               ( ndmreset_n          ),
    .boot_addr_i          ( ariane_soc::ROMBase ), // start fetching from ROM
    .core_id_i            ( '0                  ),
    .cluster_id_i         ( '0                  ),
    .irq_i                ( irq                 ),
    .ipi_i                ( ipi                 ),
    .time_irq_i           ( timer_irq           ),
    .debug_req_i          ( debug_req_irq       ),
    .data_if              ( slave_slice[2]      ),
    .bypass_if            ( slave_slice[1]      ),
    .instr_if             ( slave_slice[0]      )
);

// ---------------
// CLINT
// ---------------
// divide clock by two
always_ff @(posedge clk or negedge ndmreset_n) begin
  if (~ndmreset_n) begin
    rtc <= 0;
  end else begin
    rtc <= rtc ^ 1'b1;
  end
end

clint #(
    .AXI_ADDR_WIDTH ( AxiAddrWidth     ),
    .AXI_DATA_WIDTH ( AxiDataWidth     ),
    .AXI_ID_WIDTH   ( AxiIdWidthSlaves ),
    .NR_CORES       ( 1                )
) i_clint (
    .clk_i       ( clk                       ),
    .rst_ni      ( ndmreset_n                ),
    .slave       ( master[ariane_soc::CLINT] ),
    .rtc_i       ( rtc                       ),
    .timer_irq_o ( timer_irq                 ),
    .ipi_o       ( ipi                       )
);

// ---------------
// ROM
// ---------------
axi2mem #(
    .AXI_ID_WIDTH   ( AxiIdWidthSlaves ),
    .AXI_ADDR_WIDTH ( AxiAddrWidth     ),
    .AXI_DATA_WIDTH ( AxiDataWidth     ),
    .AXI_USER_WIDTH ( AxiUserWidth     )
) i_axi2rom (
    .clk_i  ( clk                     ),
    .rst_ni ( ndmreset_n              ),
    .slave  ( master[ariane_soc::ROM] ),
    .req_o  ( rom_req                 ),
    .we_o   (                         ),
    .addr_o ( rom_addr                ),
    .be_o   (                         ),
    .data_o (                         ),
    .data_i ( rom_rdata               )
);

bootrom i_bootrom (
    .clk_i      ( clk       ),
    .req_i      ( rom_req   ),
    .addr_i     ( rom_addr  ),
    .rdata_o    ( rom_rdata )
);

// ---------------
// Peripherals
// ---------------
ariane_peripherals #(
    .AxiAddrWidth ( AxiAddrWidth ),
    .AxiDataWidth ( AxiDataWidth ),
    `ifdef GENESYSII
    .InclSPI      ( 1'b1         ),
    `elsif VCU118
    .InclSPI      ( 1'b0         ),
    `endif
    .DummyUART    ( 1'b0         )
) i_ariane_peripherals (
    .clk_i           ( clk                      ),
    .rst_ni          ( ndmreset_n               ),
    .plic            ( master[ariane_soc::PLIC] ),
    .uart            ( master[ariane_soc::UART] ),
    .spi             ( master[ariane_soc::SPI]  ),
    .irq_o           ( irq                      ),
    .rx_i            ( rx                       ),
    .tx_o            ( tx                       ),
    .spi_clk_o       ( spi_clk_o                ),
    .spi_mosi        ( spi_mosi                 ),
    .spi_miso        ( spi_miso                 ),
    .spi_ss          ( spi_ss                   )
);

// ---------------------
// Board peripherals
// ---------------------
// ---------------
// DDR
// ---------------
logic [3:0]  s_axi_awid;
logic [63:0] s_axi_awaddr;
logic [7:0]  s_axi_awlen;
logic [2:0]  s_axi_awsize;
logic [1:0]  s_axi_awburst;
logic [0:0]  s_axi_awlock;
logic [3:0]  s_axi_awcache;
logic [2:0]  s_axi_awprot;
logic [3:0]  s_axi_awregion;
logic [3:0]  s_axi_awqos;
logic        s_axi_awvalid;
logic        s_axi_awready;
logic [63:0] s_axi_wdata;
logic [7:0]  s_axi_wstrb;
logic        s_axi_wlast;
logic        s_axi_wvalid;
logic        s_axi_wready;
logic [3:0]  s_axi_bid;
logic [1:0]  s_axi_bresp;
logic        s_axi_bvalid;
logic        s_axi_bready;
logic [3:0]  s_axi_arid;
logic [63:0] s_axi_araddr;
logic [7:0]  s_axi_arlen;
logic [2:0]  s_axi_arsize;
logic [1:0]  s_axi_arburst;
logic [0:0]  s_axi_arlock;
logic [3:0]  s_axi_arcache;
logic [2:0]  s_axi_arprot;
logic [3:0]  s_axi_arregion;
logic [3:0]  s_axi_arqos;
logic        s_axi_arvalid;
logic        s_axi_arready;
logic [3:0]  s_axi_rid;
logic [63:0] s_axi_rdata;
logic [1:0]  s_axi_rresp;
logic        s_axi_rlast;
logic        s_axi_rvalid;
logic        s_axi_rready;

assign master[ariane_soc::DRAM].r_user = '0;
assign master[ariane_soc::DRAM].b_user = '0;

axi_clock_converter_0 axi_clock_converter (
  .s_axi_aclk     ( clk                                ),
  .s_axi_aresetn  ( ndmreset_n                         ),
  .s_axi_awid     ( master[ariane_soc::DRAM].aw_id     ),
  .s_axi_awaddr   ( master[ariane_soc::DRAM].aw_addr   ),
  .s_axi_awlen    ( master[ariane_soc::DRAM].aw_len    ),
  .s_axi_awsize   ( master[ariane_soc::DRAM].aw_size   ),
  .s_axi_awburst  ( master[ariane_soc::DRAM].aw_burst  ),
  .s_axi_awlock   ( master[ariane_soc::DRAM].aw_lock   ),
  .s_axi_awcache  ( master[ariane_soc::DRAM].aw_cache  ),
  .s_axi_awprot   ( master[ariane_soc::DRAM].aw_prot   ),
  .s_axi_awregion ( master[ariane_soc::DRAM].aw_region ),
  .s_axi_awqos    ( master[ariane_soc::DRAM].aw_qos    ),
  .s_axi_awvalid  ( master[ariane_soc::DRAM].aw_valid  ),
  .s_axi_awready  ( master[ariane_soc::DRAM].aw_ready  ),
  .s_axi_wdata    ( master[ariane_soc::DRAM].w_data    ),
  .s_axi_wstrb    ( master[ariane_soc::DRAM].w_strb    ),
  .s_axi_wlast    ( master[ariane_soc::DRAM].w_last    ),
  .s_axi_wvalid   ( master[ariane_soc::DRAM].w_valid   ),
  .s_axi_wready   ( master[ariane_soc::DRAM].w_ready   ),
  .s_axi_bid      ( master[ariane_soc::DRAM].b_id      ),
  .s_axi_bresp    ( master[ariane_soc::DRAM].b_resp    ),
  .s_axi_bvalid   ( master[ariane_soc::DRAM].b_valid   ),
  .s_axi_bready   ( master[ariane_soc::DRAM].b_ready   ),
  .s_axi_arid     ( master[ariane_soc::DRAM].ar_id     ),
  .s_axi_araddr   ( master[ariane_soc::DRAM].ar_addr   ),
  .s_axi_arlen    ( master[ariane_soc::DRAM].ar_len    ),
  .s_axi_arsize   ( master[ariane_soc::DRAM].ar_size   ),
  .s_axi_arburst  ( master[ariane_soc::DRAM].ar_burst  ),
  .s_axi_arlock   ( master[ariane_soc::DRAM].ar_lock   ),
  .s_axi_arcache  ( master[ariane_soc::DRAM].ar_cache  ),
  .s_axi_arprot   ( master[ariane_soc::DRAM].ar_prot   ),
  .s_axi_arregion ( master[ariane_soc::DRAM].ar_region ),
  .s_axi_arqos    ( master[ariane_soc::DRAM].ar_qos    ),
  .s_axi_arvalid  ( master[ariane_soc::DRAM].ar_valid  ),
  .s_axi_arready  ( master[ariane_soc::DRAM].ar_ready  ),
  .s_axi_rid      ( master[ariane_soc::DRAM].r_id      ),
  .s_axi_rdata    ( master[ariane_soc::DRAM].r_data    ),
  .s_axi_rresp    ( master[ariane_soc::DRAM].r_resp    ),
  .s_axi_rlast    ( master[ariane_soc::DRAM].r_last    ),
  .s_axi_rvalid   ( master[ariane_soc::DRAM].r_valid   ),
  .s_axi_rready   ( master[ariane_soc::DRAM].r_ready   ),
  // to size converter
  .m_axi_aclk     ( ddr_clock_out                      ),
  .m_axi_aresetn  ( ndmreset_n                         ),
  .m_axi_awid     ( s_axi_awid                         ),
  .m_axi_awaddr   ( s_axi_awaddr                       ),
  .m_axi_awlen    ( s_axi_awlen                        ),
  .m_axi_awsize   ( s_axi_awsize                       ),
  .m_axi_awburst  ( s_axi_awburst                      ),
  .m_axi_awlock   ( s_axi_awlock                       ),
  .m_axi_awcache  ( s_axi_awcache                      ),
  .m_axi_awprot   ( s_axi_awprot                       ),
  .m_axi_awregion ( s_axi_awregion                     ),
  .m_axi_awqos    ( s_axi_awqos                        ),
  .m_axi_awvalid  ( s_axi_awvalid                      ),
  .m_axi_awready  ( s_axi_awready                      ),
  .m_axi_wdata    ( s_axi_wdata                        ),
  .m_axi_wstrb    ( s_axi_wstrb                        ),
  .m_axi_wlast    ( s_axi_wlast                        ),
  .m_axi_wvalid   ( s_axi_wvalid                       ),
  .m_axi_wready   ( s_axi_wready                       ),
  .m_axi_bid      ( s_axi_bid                          ),
  .m_axi_bresp    ( s_axi_bresp                        ),
  .m_axi_bvalid   ( s_axi_bvalid                       ),
  .m_axi_bready   ( s_axi_bready                       ),
  .m_axi_arid     ( s_axi_arid                         ),
  .m_axi_araddr   ( s_axi_araddr                       ),
  .m_axi_arlen    ( s_axi_arlen                        ),
  .m_axi_arsize   ( s_axi_arsize                       ),
  .m_axi_arburst  ( s_axi_arburst                      ),
  .m_axi_arlock   ( s_axi_arlock                       ),
  .m_axi_arcache  ( s_axi_arcache                      ),
  .m_axi_arprot   ( s_axi_arprot                       ),
  .m_axi_arregion ( s_axi_arregion                     ),
  .m_axi_arqos    ( s_axi_arqos                        ),
  .m_axi_arvalid  ( s_axi_arvalid                      ),
  .m_axi_arready  ( s_axi_arready                      ),
  .m_axi_rid      ( s_axi_rid                          ),
  .m_axi_rdata    ( s_axi_rdata                        ),
  .m_axi_rresp    ( s_axi_rresp                        ),
  .m_axi_rlast    ( s_axi_rlast                        ),
  .m_axi_rvalid   ( s_axi_rvalid                       ),
  .m_axi_rready   ( s_axi_rready                       )
);

clk_wiz_0 i_clk_gen (
  .clk_out1 ( clk           ),
  .reset    ( cpu_reset     ),
  .locked   (               ), // keep open
  .clk_in1  ( ddr_clock_out )
);

`ifdef INCL_SRAM
  logic                       req;
  logic                       we;
  logic [AxiAddrWidth-1:0]    addr;
  logic [AxiDataWidth/8-1:0]  be;
  logic [AxiDataWidth-1:0]    wdata;
  logic [AxiDataWidth-1:0]    rdata;

  axi2mem #(
      .AXI_ID_WIDTH   ( AxiIdWidthSlaves ),
      .AXI_ADDR_WIDTH ( AxiAddrWidth     ),
      .AXI_DATA_WIDTH ( AxiDataWidth     ),
      .AXI_USER_WIDTH ( AxiUserWidth     )
  ) i_axi2mem (
      .clk_i  ( clk                      ),
      .rst_ni ( ndmreset_n               ),
      .slave  ( master[ariane_soc::DRAM] ),
      .req_o  ( req                      ),
      .we_o   ( we                       ),
      .addr_o ( addr                     ),
      .be_o   ( be                       ),
      .data_o ( wdata                    ),
      .data_i ( rdata                    )
  );

  // sram #(
  //     .DATA_WIDTH ( AxiDataWidth ),
  //     .NUM_WORDS  ( NumWords     )
  // ) i_sram (
  //     .clk_i      ( clk                                                                    ),
  //     .rst_ni     ( rst_ni                                                                 ),
  //     .req_i      ( req                                                                    ),
  //     .we_i       ( we                                                                     ),
  //     .addr_i     ( addr[$clog2(NumWords)-1+$clog2(AxiDataWidth/8):$clog2(AxiDataWidth/8)] ),
  //     .wdata_i    ( wdata                                                                  ),
  //     .be_i       ( be                                                                     ),
  //     .rdata_o    ( rdata                                                                  )
  // );
  xpm_memory_spram #(
    .ADDR_WIDTH_A        ( $clog2(NumWords) ),
    .AUTO_SLEEP_TIME     ( 0                ),
    .BYTE_WRITE_WIDTH_A  ( 8                ),
    .ECC_MODE            ( "no_ecc"         ),
    .MEMORY_OPTIMIZATION ( "true"           ),
    .MEMORY_PRIMITIVE    ( "auto"           ),
    .MEMORY_SIZE         ( NumWords * 64    ),
    .MESSAGE_CONTROL     ( 0                ),
    .READ_DATA_WIDTH_A   ( 64               ),
    .READ_LATENCY_A      ( 1                ),
    .USE_MEM_INIT        ( 0                ),
    .WAKEUP_TIME         ( "disable_sleep"  ),
    .WRITE_DATA_WIDTH_A  ( 64               ),
    .WRITE_MODE_A        ( "read_first"     )
  ) xpm_memory_spram_inst (
    .dbiterra       (                                                                        ),
    .douta          ( rdata                                                                  ),
    .sbiterra       (                                                                        ),
    .addra          ( addr[$clog2(NumWords)-1+$clog2(AxiDataWidth/8):$clog2(AxiDataWidth/8)] ),
    .clka           ( clk                                                                    ),
    .dina           ( wdata                                                                  ),
    .ena            ( req                                                                    ),
    .injectdbiterra ( '0                                                                     ),
    .injectsbiterra ( '0                                                                     ),
    .regcea         ( 1'b1                                                                   ),
    .rsta           ( rst                                                                    ),
    .sleep          ( 1'b0                                                                   ),
    .wea            ( we                                                                     )
  );
`endif

`ifdef GENESYSII
fan_ctrl i_fan_ctrl (
    .clk_i         ( clk        ),
    .rst_ni        ( ndmreset_n ),
    .pwm_setting_i ( sw[3:0]    ),
    .fan_pwm_o     ( fan_pwm    )
);

ariane_leds i_ariane_leds (
  .clk_i          ( clk          ),
  .rst_ni         ( rst_n        ),
  .led_o          ( led          ),
  .pc_asserted_i  ( pc_asserted  ),
  .dmactive_i     ( dmactive     ),
  .commit_valid_i ( '0           )
);

mig_7series_0 i_ddr (
    .sys_clk_p,
    .sys_clk_n,
    .ddr3_dq,
    .ddr3_dqs_n,
    .ddr3_dqs_p,
    .ddr3_addr,
    .ddr3_ba,
    .ddr3_ras_n,
    .ddr3_cas_n,
    .ddr3_we_n,
    .ddr3_reset_n,
    .ddr3_ck_p,
    .ddr3_ck_n,
    .ddr3_cke,
    .ddr3_cs_n,
    .ddr3_dm,
    .ddr3_odt,
    .mmcm_locked     (                ), // keep open
    .app_sr_req      ( '0             ),
    .app_ref_req     ( '0             ),
    .app_zq_req      ( '0             ),
    .app_sr_active   (                ), // keep open
    .app_ref_ack     (                ), // keep open
    .app_zq_ack      (                ), // keep open
    .ui_clk          ( ddr_clock_out  ),
    .ui_clk_sync_rst ( ddr_sync_reset ),
    .aresetn         ( ndmreset_n     ),
    .s_axi_awid,
    .s_axi_awaddr    ( s_axi_awaddr[29:0] ),
    .s_axi_awlen,
    .s_axi_awsize,
    .s_axi_awburst,
    .s_axi_awlock,
    .s_axi_awcache,
    .s_axi_awprot,
    .s_axi_awqos,
    .s_axi_awvalid,
    .s_axi_awready,
    .s_axi_wdata,
    .s_axi_wstrb,
    .s_axi_wlast,
    .s_axi_wvalid,
    .s_axi_wready,
    .s_axi_bready,
    .s_axi_bid,
    .s_axi_bresp,
    .s_axi_bvalid,
    .s_axi_arid,
    .s_axi_araddr     ( s_axi_araddr[29:0] ),
    .s_axi_arlen,
    .s_axi_arsize,
    .s_axi_arburst,
    .s_axi_arlock,
    .s_axi_arcache,
    .s_axi_arprot,
    .s_axi_arqos,
    .s_axi_arvalid,
    .s_axi_arready,
    .s_axi_rready,
    .s_axi_rid,
    .s_axi_rdata,
    .s_axi_rresp,
    .s_axi_rlast,
    .s_axi_rvalid,
    .init_calib_complete (            ), // keep open
    .device_temp         (            ), // keep open
    .sys_rst             ( cpu_resetn )
);
`elsif VCU118

  logic [63:0]  dram_dwidth_axi_awaddr;
  logic [7:0]   dram_dwidth_axi_awlen;
  logic [2:0]   dram_dwidth_axi_awsize;
  logic [1:0]   dram_dwidth_axi_awburst;
  logic [0:0]   dram_dwidth_axi_awlock;
  logic [3:0]   dram_dwidth_axi_awcache;
  logic [2:0]   dram_dwidth_axi_awprot;
  logic [3:0]   dram_dwidth_axi_awqos;
  logic         dram_dwidth_axi_awvalid;
  logic         dram_dwidth_axi_awready;
  logic [511:0] dram_dwidth_axi_wdata;
  logic [63:0]  dram_dwidth_axi_wstrb;
  logic         dram_dwidth_axi_wlast;
  logic         dram_dwidth_axi_wvalid;
  logic         dram_dwidth_axi_wready;
  logic         dram_dwidth_axi_bready;
  logic [1:0]   dram_dwidth_axi_bresp;
  logic         dram_dwidth_axi_bvalid;
  logic [63:0]  dram_dwidth_axi_araddr;
  logic [7:0]   dram_dwidth_axi_arlen;
  logic [2:0]   dram_dwidth_axi_arsize;
  logic [1:0]   dram_dwidth_axi_arburst;
  logic [0:0]   dram_dwidth_axi_arlock;
  logic [3:0]   dram_dwidth_axi_arcache;
  logic [2:0]   dram_dwidth_axi_arprot;
  logic [3:0]   dram_dwidth_axi_arqos;
  logic         dram_dwidth_axi_arvalid;
  logic         dram_dwidth_axi_arready;
  logic         dram_dwidth_axi_rready;
  logic         dram_dwidth_axi_rlast;
  logic         dram_dwidth_axi_rvalid;
  logic [1:0]   dram_dwidth_axi_rresp;
  logic [511:0] dram_dwidth_axi_rdata;

axi_dwidth_converter_512_64 i_axi_dwidth_converter_512_64 (
  .s_axi_aclk     ( ddr_clock_out            ),
  .s_axi_aresetn  ( rst_n                    ),

  .s_axi_awid     ( s_axi_awid               ),
  .s_axi_awaddr   ( s_axi_awaddr             ),
  .s_axi_awlen    ( s_axi_awlen              ),
  .s_axi_awsize   ( s_axi_awsize             ),
  .s_axi_awburst  ( s_axi_awburst            ),
  .s_axi_awlock   ( s_axi_awlock             ),
  .s_axi_awcache  ( s_axi_awcache            ),
  .s_axi_awprot   ( s_axi_awprot             ),
  .s_axi_awregion ( '0                       ),
  .s_axi_awqos    ( s_axi_awqos              ),
  .s_axi_awvalid  ( s_axi_awvalid            ),
  .s_axi_awready  ( s_axi_awready            ),
  .s_axi_wdata    ( s_axi_wdata              ),
  .s_axi_wstrb    ( s_axi_wstrb              ),
  .s_axi_wlast    ( s_axi_wlast              ),
  .s_axi_wvalid   ( s_axi_wvalid             ),
  .s_axi_wready   ( s_axi_wready             ),
  .s_axi_bid      ( s_axi_bid                ),
  .s_axi_bresp    ( s_axi_bresp              ),
  .s_axi_bvalid   ( s_axi_bvalid             ),
  .s_axi_bready   ( s_axi_bready             ),
  .s_axi_arid     ( s_axi_arid               ),
  .s_axi_araddr   ( s_axi_araddr             ),
  .s_axi_arlen    ( s_axi_arlen              ),
  .s_axi_arsize   ( s_axi_arsize             ),
  .s_axi_arburst  ( s_axi_arburst            ),
  .s_axi_arlock   ( s_axi_arlock             ),
  .s_axi_arcache  ( s_axi_arcache            ),
  .s_axi_arprot   ( s_axi_arprot             ),
  .s_axi_arregion ( '0                       ),
  .s_axi_arqos    ( s_axi_arqos              ),
  .s_axi_arvalid  ( s_axi_arvalid            ),
  .s_axi_arready  ( s_axi_arready            ),
  .s_axi_rid      ( s_axi_rid                ),
  .s_axi_rdata    ( s_axi_rdata              ),
  .s_axi_rresp    ( s_axi_rresp              ),
  .s_axi_rlast    ( s_axi_rlast              ),
  .s_axi_rvalid   ( s_axi_rvalid             ),
  .s_axi_rready   ( s_axi_rready             ),

  .m_axi_awaddr   ( dram_dwidth_axi_awaddr   ),
  .m_axi_awlen    ( dram_dwidth_axi_awlen    ),
  .m_axi_awsize   ( dram_dwidth_axi_awsize   ),
  .m_axi_awburst  ( dram_dwidth_axi_awburst  ),
  .m_axi_awlock   ( dram_dwidth_axi_awlock   ),
  .m_axi_awcache  ( dram_dwidth_axi_awcache  ),
  .m_axi_awprot   ( dram_dwidth_axi_awprot   ),
  .m_axi_awregion (                          ), // left open
  .m_axi_awqos    ( dram_dwidth_axi_awqos    ),
  .m_axi_awvalid  ( dram_dwidth_axi_awvalid  ),
  .m_axi_awready  ( dram_dwidth_axi_awready  ),
  .m_axi_wdata    ( dram_dwidth_axi_wdata    ),
  .m_axi_wstrb    ( dram_dwidth_axi_wstrb    ),
  .m_axi_wlast    ( dram_dwidth_axi_wlast    ),
  .m_axi_wvalid   ( dram_dwidth_axi_wvalid   ),
  .m_axi_wready   ( dram_dwidth_axi_wready   ),
  .m_axi_bresp    ( dram_dwidth_axi_bresp    ),
  .m_axi_bvalid   ( dram_dwidth_axi_bvalid   ),
  .m_axi_bready   ( dram_dwidth_axi_bready   ),
  .m_axi_araddr   ( dram_dwidth_axi_araddr   ),
  .m_axi_arlen    ( dram_dwidth_axi_arlen    ),
  .m_axi_arsize   ( dram_dwidth_axi_arsize   ),
  .m_axi_arburst  ( dram_dwidth_axi_arburst  ),
  .m_axi_arlock   ( dram_dwidth_axi_arlock   ),
  .m_axi_arcache  ( dram_dwidth_axi_arcache  ),
  .m_axi_arprot   ( dram_dwidth_axi_arprot   ),
  .m_axi_arregion (                          ),
  .m_axi_arqos    ( dram_dwidth_axi_arqos    ),
  .m_axi_arvalid  ( dram_dwidth_axi_arvalid  ),
  .m_axi_arready  ( dram_dwidth_axi_arready  ),
  .m_axi_rdata    ( dram_dwidth_axi_rdata    ),
  .m_axi_rresp    ( dram_dwidth_axi_rresp    ),
  .m_axi_rlast    ( dram_dwidth_axi_rlast    ),
  .m_axi_rvalid   ( dram_dwidth_axi_rvalid   ),
  .m_axi_rready   ( dram_dwidth_axi_rready   )
);

  ddr4_0 i_ddr (
    .c0_init_calib_complete (                              ),
    .dbg_clk                (                              ),
    .c0_sys_clk_p           ( c0_sys_clk_p                 ),
    .c0_sys_clk_n           ( c0_sys_clk_n                 ),
    .dbg_bus                (                              ),
    .c0_ddr4_adr            ( c0_ddr4_adr                  ),
    .c0_ddr4_ba             ( c0_ddr4_ba                   ),
    .c0_ddr4_cke            ( c0_ddr4_cke                  ),
    .c0_ddr4_cs_n           ( c0_ddr4_cs_n                 ),
    .c0_ddr4_dm_dbi_n       ( c0_ddr4_dm_dbi_n             ),
    .c0_ddr4_dq             ( c0_ddr4_dq                   ),
    .c0_ddr4_dqs_c          ( c0_ddr4_dqs_c                ),
    .c0_ddr4_dqs_t          ( c0_ddr4_dqs_t                ),
    .c0_ddr4_odt            ( c0_ddr4_odt                  ),
    .c0_ddr4_bg             ( c0_ddr4_bg                   ),
    .c0_ddr4_reset_n        ( c0_ddr4_reset_n              ),
    .c0_ddr4_act_n          ( c0_ddr4_act_n                ),
    .c0_ddr4_ck_c           ( c0_ddr4_ck_c                 ),
    .c0_ddr4_ck_t           ( c0_ddr4_ck_t                 ),
    .c0_ddr4_ui_clk         ( ddr_clock_out                ),
    .c0_ddr4_ui_clk_sync_rst( ddr_sync_reset               ),
    .c0_ddr4_aresetn        ( ndmreset_n                   ),
    .c0_ddr4_s_axi_awid     ( '0                           ),
    .c0_ddr4_s_axi_awaddr   ( dram_dwidth_axi_awaddr[30:0] ),
    .c0_ddr4_s_axi_awlen    ( dram_dwidth_axi_awlen        ),
    .c0_ddr4_s_axi_awsize   ( dram_dwidth_axi_awsize       ),
    .c0_ddr4_s_axi_awburst  ( dram_dwidth_axi_awburst      ),
    .c0_ddr4_s_axi_awlock   ( dram_dwidth_axi_awlock       ),
    .c0_ddr4_s_axi_awcache  ( dram_dwidth_axi_awcache      ),
    .c0_ddr4_s_axi_awprot   ( dram_dwidth_axi_awprot       ),
    .c0_ddr4_s_axi_awqos    ( dram_dwidth_axi_awqos        ),
    .c0_ddr4_s_axi_awvalid  ( dram_dwidth_axi_awvalid      ),
    .c0_ddr4_s_axi_awready  ( dram_dwidth_axi_awready      ),
    .c0_ddr4_s_axi_wdata    ( dram_dwidth_axi_wdata        ),
    .c0_ddr4_s_axi_wstrb    ( dram_dwidth_axi_wstrb        ),
    .c0_ddr4_s_axi_wlast    ( dram_dwidth_axi_wlast        ),
    .c0_ddr4_s_axi_wvalid   ( dram_dwidth_axi_wvalid       ),
    .c0_ddr4_s_axi_wready   ( dram_dwidth_axi_wready       ),
    .c0_ddr4_s_axi_bready   ( dram_dwidth_axi_bready       ),
    .c0_ddr4_s_axi_bid      (                              ),
    .c0_ddr4_s_axi_bresp    ( dram_dwidth_axi_bresp        ),
    .c0_ddr4_s_axi_bvalid   ( dram_dwidth_axi_bvalid       ),
    .c0_ddr4_s_axi_arid     ( '0                           ),
    .c0_ddr4_s_axi_araddr   ( dram_dwidth_axi_araddr[30:0] ),
    .c0_ddr4_s_axi_arlen    ( dram_dwidth_axi_arlen        ),
    .c0_ddr4_s_axi_arsize   ( dram_dwidth_axi_arsize       ),
    .c0_ddr4_s_axi_arburst  ( dram_dwidth_axi_arburst      ),
    .c0_ddr4_s_axi_arlock   ( dram_dwidth_axi_arlock       ),
    .c0_ddr4_s_axi_arcache  ( dram_dwidth_axi_arcache      ),
    .c0_ddr4_s_axi_arprot   ( dram_dwidth_axi_arprot       ),
    .c0_ddr4_s_axi_arqos    ( dram_dwidth_axi_arqos        ),
    .c0_ddr4_s_axi_arvalid  ( dram_dwidth_axi_arvalid      ),
    .c0_ddr4_s_axi_arready  ( dram_dwidth_axi_arready      ),
    .c0_ddr4_s_axi_rready   ( dram_dwidth_axi_rready       ),
    .c0_ddr4_s_axi_rlast    ( dram_dwidth_axi_rlast        ),
    .c0_ddr4_s_axi_rvalid   ( dram_dwidth_axi_rvalid       ),
    .c0_ddr4_s_axi_rresp    ( dram_dwidth_axi_rresp        ),
    .c0_ddr4_s_axi_rid      (                              ),
    .c0_ddr4_s_axi_rdata    ( dram_dwidth_axi_rdata        ),
    .sys_rst                ( cpu_reset                    )
  );


  logic pcie_ref_clk;
  logic pcie_ref_clk_gt;

  logic pcie_axi_clk;
  logic pcie_axi_rstn;

  logic         pcie_axi_awready;
  logic         pcie_axi_wready;
  logic [3:0]   pcie_axi_bid;
  logic [1:0]   pcie_axi_bresp;
  logic         pcie_axi_bvalid;
  logic         pcie_axi_arready;
  logic [3:0]   pcie_axi_rid;
  logic [255:0] pcie_axi_rdata;
  logic [1:0]   pcie_axi_rresp;
  logic         pcie_axi_rlast;
  logic         pcie_axi_rvalid;
  logic [3:0]   pcie_axi_awid;
  logic [63:0]  pcie_axi_awaddr;
  logic [7:0]   pcie_axi_awlen;
  logic [2:0]   pcie_axi_awsize;
  logic [1:0]   pcie_axi_awburst;
  logic [2:0]   pcie_axi_awprot;
  logic         pcie_axi_awvalid;
  logic         pcie_axi_awlock;
  logic [3:0]   pcie_axi_awcache;
  logic [255:0] pcie_axi_wdata;
  logic [31:0]  pcie_axi_wstrb;
  logic         pcie_axi_wlast;
  logic         pcie_axi_wvalid;
  logic         pcie_axi_bready;
  logic [3:0]   pcie_axi_arid;
  logic [63:0]  pcie_axi_araddr;
  logic [7:0]   pcie_axi_arlen;
  logic [2:0]   pcie_axi_arsize;
  logic [1:0]   pcie_axi_arburst;
  logic [2:0]   pcie_axi_arprot;
  logic         pcie_axi_arvalid;
  logic         pcie_axi_arlock;
  logic [3:0]   pcie_axi_arcache;
  logic         pcie_axi_rready;

  logic [63:0]  pcie_dwidth_axi_awaddr;
  logic [7:0]   pcie_dwidth_axi_awlen;
  logic [2:0]   pcie_dwidth_axi_awsize;
  logic [1:0]   pcie_dwidth_axi_awburst;
  logic [0:0]   pcie_dwidth_axi_awlock;
  logic [3:0]   pcie_dwidth_axi_awcache;
  logic [2:0]   pcie_dwidth_axi_awprot;
  logic [3:0]   pcie_dwidth_axi_awregion;
  logic [3:0]   pcie_dwidth_axi_awqos;
  logic         pcie_dwidth_axi_awvalid;
  logic         pcie_dwidth_axi_awready;
  logic [63:0]  pcie_dwidth_axi_wdata;
  logic [7:0]   pcie_dwidth_axi_wstrb;
  logic         pcie_dwidth_axi_wlast;
  logic         pcie_dwidth_axi_wvalid;
  logic         pcie_dwidth_axi_wready;
  logic [1:0]   pcie_dwidth_axi_bresp;
  logic         pcie_dwidth_axi_bvalid;
  logic         pcie_dwidth_axi_bready;
  logic [63:0]  pcie_dwidth_axi_araddr;
  logic [7:0]   pcie_dwidth_axi_arlen;
  logic [2:0]   pcie_dwidth_axi_arsize;
  logic [1:0]   pcie_dwidth_axi_arburst;
  logic [0:0]   pcie_dwidth_axi_arlock;
  logic [3:0]   pcie_dwidth_axi_arcache;
  logic [2:0]   pcie_dwidth_axi_arprot;
  logic [3:0]   pcie_dwidth_axi_arregion;
  logic [3:0]   pcie_dwidth_axi_arqos;
  logic         pcie_dwidth_axi_arvalid;
  logic         pcie_dwidth_axi_arready;
  logic [63:0]  pcie_dwidth_axi_rdata;
  logic [1:0]   pcie_dwidth_axi_rresp;
  logic         pcie_dwidth_axi_rlast;
  logic         pcie_dwidth_axi_rvalid;
  logic         pcie_dwidth_axi_rready;

  // PCIe Reset
  logic sys_rst_n_c;
  IBUF sys_reset_n_ibuf (.O(sys_rst_n_c), .I(sys_rst_n));

  IBUFDS_GTE4 #(
    .REFCLK_HROW_CK_SEL ( 2'b00 )
  ) IBUFDS_GTE4_inst (
    .O     ( pcie_ref_clk_gt ),
    .ODIV2 ( pcie_ref_clk    ),
    .CEB   ( 1'b0            ),
    .I     ( sys_clk_p       ),
    .IB    ( sys_clk_n       )
  );

  // 250 MHz AXI
  xdma_0 i_xdma (
    .sys_clk                  ( pcie_ref_clk     ),
    .sys_clk_gt               ( pcie_ref_clk_gt  ),
    .sys_rst_n                ( sys_rst_n_c      ),
    .user_lnk_up              (                  ),

    // Tx
    .pci_exp_txp              ( pci_exp_txp      ),
    .pci_exp_txn              ( pci_exp_txn      ),
    // Rx
    .pci_exp_rxp              ( pci_exp_rxp      ),
    .pci_exp_rxn              ( pci_exp_rxn      ),
    .usr_irq_req              ( 1'b0             ),
    .usr_irq_ack              (                  ),
    .msi_enable               (                  ),
    .msi_vector_width         (                  ),
    .axi_aclk                 ( pcie_axi_clk     ),
    .axi_aresetn              ( pcie_axi_rstn    ),
    .m_axi_awready            ( pcie_axi_awready ),
    .m_axi_wready             ( pcie_axi_wready  ),
    .m_axi_bid                ( pcie_axi_bid     ),
    .m_axi_bresp              ( pcie_axi_bresp   ),
    .m_axi_bvalid             ( pcie_axi_bvalid  ),
    .m_axi_arready            ( pcie_axi_arready ),
    .m_axi_rid                ( pcie_axi_rid     ),
    .m_axi_rdata              ( pcie_axi_rdata   ),
    .m_axi_rresp              ( pcie_axi_rresp   ),
    .m_axi_rlast              ( pcie_axi_rlast   ),
    .m_axi_rvalid             ( pcie_axi_rvalid  ),
    .m_axi_awid               ( pcie_axi_awid    ),
    .m_axi_awaddr             ( pcie_axi_awaddr  ),
    .m_axi_awlen              ( pcie_axi_awlen   ),
    .m_axi_awsize             ( pcie_axi_awsize  ),
    .m_axi_awburst            ( pcie_axi_awburst ),
    .m_axi_awprot             ( pcie_axi_awprot  ),
    .m_axi_awvalid            ( pcie_axi_awvalid ),
    .m_axi_awlock             ( pcie_axi_awlock  ),
    .m_axi_awcache            ( pcie_axi_awcache ),
    .m_axi_wdata              ( pcie_axi_wdata   ),
    .m_axi_wstrb              ( pcie_axi_wstrb   ),
    .m_axi_wlast              ( pcie_axi_wlast   ),
    .m_axi_wvalid             ( pcie_axi_wvalid  ),
    .m_axi_bready             ( pcie_axi_bready  ),
    .m_axi_arid               ( pcie_axi_arid    ),
    .m_axi_araddr             ( pcie_axi_araddr  ),
    .m_axi_arlen              ( pcie_axi_arlen   ),
    .m_axi_arsize             ( pcie_axi_arsize  ),
    .m_axi_arburst            ( pcie_axi_arburst ),
    .m_axi_arprot             ( pcie_axi_arprot  ),
    .m_axi_arvalid            ( pcie_axi_arvalid ),
    .m_axi_arlock             ( pcie_axi_arlock  ),
    .m_axi_arcache            ( pcie_axi_arcache ),
    .m_axi_rready             ( pcie_axi_rready  ),

    .cfg_mgmt_addr            ( '0               ),
    .cfg_mgmt_write           ( '0               ),
    .cfg_mgmt_write_data      ( '0               ),
    .cfg_mgmt_byte_enable     ( '0               ),
    .cfg_mgmt_read            ( '0               ),
    .cfg_mgmt_read_data       (                  ),
    .cfg_mgmt_read_write_done (                  )
  );

  axi_dwidth_converter_256_64 i_axi_dwidth_converter_256_64 (
    .s_axi_aclk     ( pcie_axi_clk             ),
    .s_axi_aresetn  ( pcie_axi_rstn            ),
    .s_axi_awid     ( pcie_axi_awid            ),
    .s_axi_awaddr   ( pcie_axi_awaddr          ),
    .s_axi_awlen    ( pcie_axi_awlen           ),
    .s_axi_awsize   ( pcie_axi_awsize          ),
    .s_axi_awburst  ( pcie_axi_awburst         ),
    .s_axi_awlock   ( pcie_axi_awlock          ),
    .s_axi_awcache  ( pcie_axi_awcache         ),
    .s_axi_awprot   ( pcie_axi_awprot          ),
    .s_axi_awregion ( '0                       ),
    .s_axi_awqos    ( '0                       ),
    .s_axi_awvalid  ( pcie_axi_awvalid         ),
    .s_axi_awready  ( pcie_axi_awready         ),
    .s_axi_wdata    ( pcie_axi_wdata           ),
    .s_axi_wstrb    ( pcie_axi_wstrb           ),
    .s_axi_wlast    ( pcie_axi_wlast           ),
    .s_axi_wvalid   ( pcie_axi_wvalid          ),
    .s_axi_wready   ( pcie_axi_wready          ),
    .s_axi_bid      ( pcie_axi_bid             ),
    .s_axi_bresp    ( pcie_axi_rresp           ),
    .s_axi_bvalid   ( pcie_axi_bvalid          ),
    .s_axi_bready   ( pcie_axi_bready          ),
    .s_axi_arid     ( pcie_axi_arid            ),
    .s_axi_araddr   ( pcie_axi_araddr          ),
    .s_axi_arlen    ( pcie_axi_arlen           ),
    .s_axi_arsize   ( pcie_axi_arsize          ),
    .s_axi_arburst  ( pcie_axi_arburst         ),
    .s_axi_arlock   ( pcie_axi_arlock          ),
    .s_axi_arcache  ( pcie_axi_arcache         ),
    .s_axi_arprot   ( pcie_axi_arprot          ),
    .s_axi_arregion ( '0                       ),
    .s_axi_arqos    ( '0                       ),
    .s_axi_arvalid  ( pcie_axi_arvalid         ),
    .s_axi_arready  ( pcie_axi_arready         ),
    .s_axi_rid      ( pcie_axi_rid             ),
    .s_axi_rdata    ( pcie_axi_rdata           ),
    .s_axi_rresp    ( pcie_axi_bresp           ),
    .s_axi_rlast    ( pcie_axi_rlast           ),
    .s_axi_rvalid   ( pcie_axi_rvalid          ),
    .s_axi_rready   ( pcie_axi_rready          ),

    .m_axi_awaddr   ( pcie_dwidth_axi_awaddr   ),
    .m_axi_awlen    ( pcie_dwidth_axi_awlen    ),
    .m_axi_awsize   ( pcie_dwidth_axi_awsize   ),
    .m_axi_awburst  ( pcie_dwidth_axi_awburst  ),
    .m_axi_awlock   ( pcie_dwidth_axi_awlock   ),
    .m_axi_awcache  ( pcie_dwidth_axi_awcache  ),
    .m_axi_awprot   ( pcie_dwidth_axi_awprot   ),
    .m_axi_awregion ( pcie_dwidth_axi_awregion ),
    .m_axi_awqos    ( pcie_dwidth_axi_awqos    ),
    .m_axi_awvalid  ( pcie_dwidth_axi_awvalid  ),
    .m_axi_awready  ( pcie_dwidth_axi_awready  ),
    .m_axi_wdata    ( pcie_dwidth_axi_wdata    ),
    .m_axi_wstrb    ( pcie_dwidth_axi_wstrb    ),
    .m_axi_wlast    ( pcie_dwidth_axi_wlast    ),
    .m_axi_wvalid   ( pcie_dwidth_axi_wvalid   ),
    .m_axi_wready   ( pcie_dwidth_axi_wready   ),
    .m_axi_bresp    ( pcie_dwidth_axi_bresp    ),
    .m_axi_bvalid   ( pcie_dwidth_axi_bvalid   ),
    .m_axi_bready   ( pcie_dwidth_axi_bready   ),
    .m_axi_araddr   ( pcie_dwidth_axi_araddr   ),
    .m_axi_arlen    ( pcie_dwidth_axi_arlen    ),
    .m_axi_arsize   ( pcie_dwidth_axi_arsize   ),
    .m_axi_arburst  ( pcie_dwidth_axi_arburst  ),
    .m_axi_arlock   ( pcie_dwidth_axi_arlock   ),
    .m_axi_arcache  ( pcie_dwidth_axi_arcache  ),
    .m_axi_arprot   ( pcie_dwidth_axi_arprot   ),
    .m_axi_arregion ( pcie_dwidth_axi_arregion ),
    .m_axi_arqos    ( pcie_dwidth_axi_arqos    ),
    .m_axi_arvalid  ( pcie_dwidth_axi_arvalid  ),
    .m_axi_arready  ( pcie_dwidth_axi_arready  ),
    .m_axi_rdata    ( pcie_dwidth_axi_rdata    ),
    .m_axi_rresp    ( pcie_dwidth_axi_rresp    ),
    .m_axi_rlast    ( pcie_dwidth_axi_rlast    ),
    .m_axi_rvalid   ( pcie_dwidth_axi_rvalid   ),
    .m_axi_rready   ( pcie_dwidth_axi_rready   )
  );


assign slave_slice[3].aw_user = '0;
assign slave_slice[3].ar_user = '0;
assign slave_slice[3].w_user = '0;

logic [3:0] slave_slice_b_id;
logic [3:0] slave_slice_r_id;

assign slave_slice[3].b_id = slave_slice_b_id[1:0];
assign slave_slice[3].r_id = slave_slice_r_id[1:0];

// PCIe Clock Converter
axi_clock_converter_0 pcie_axi_clock_converter (
  .m_axi_aclk     ( clk                      ),
  .m_axi_aresetn  ( ndmreset_n               ),
  .m_axi_awid     ( {2'b0, slave_slice[3].aw_id} ),
  .m_axi_awaddr   ( slave_slice[3].aw_addr   ),
  .m_axi_awlen    ( slave_slice[3].aw_len    ),
  .m_axi_awsize   ( slave_slice[3].aw_size   ),
  .m_axi_awburst  ( slave_slice[3].aw_burst  ),
  .m_axi_awlock   ( slave_slice[3].aw_lock   ),
  .m_axi_awcache  ( slave_slice[3].aw_cache  ),
  .m_axi_awprot   ( slave_slice[3].aw_prot   ),
  .m_axi_awregion ( slave_slice[3].aw_region ),
  .m_axi_awqos    ( slave_slice[3].aw_qos    ),
  .m_axi_awvalid  ( slave_slice[3].aw_valid  ),
  .m_axi_awready  ( slave_slice[3].aw_ready  ),
  .m_axi_wdata    ( slave_slice[3].w_data    ),
  .m_axi_wstrb    ( slave_slice[3].w_strb    ),
  .m_axi_wlast    ( slave_slice[3].w_last    ),
  .m_axi_wvalid   ( slave_slice[3].w_valid   ),
  .m_axi_wready   ( slave_slice[3].w_ready   ),
  .m_axi_bid      ( slave_slice_b_id         ),
  .m_axi_bresp    ( slave_slice[3].b_resp    ),
  .m_axi_bvalid   ( slave_slice[3].b_valid   ),
  .m_axi_bready   ( slave_slice[3].b_ready   ),
  .m_axi_arid     ( {2'b0, slave_slice[3].ar_id} ),
  .m_axi_araddr   ( slave_slice[3].ar_addr   ),
  .m_axi_arlen    ( slave_slice[3].ar_len    ),
  .m_axi_arsize   ( slave_slice[3].ar_size   ),
  .m_axi_arburst  ( slave_slice[3].ar_burst  ),
  .m_axi_arlock   ( slave_slice[3].ar_lock   ),
  .m_axi_arcache  ( slave_slice[3].ar_cache  ),
  .m_axi_arprot   ( slave_slice[3].ar_prot   ),
  .m_axi_arregion ( slave_slice[3].ar_region ),
  .m_axi_arqos    ( slave_slice[3].ar_qos    ),
  .m_axi_arvalid  ( slave_slice[3].ar_valid  ),
  .m_axi_arready  ( slave_slice[3].ar_ready  ),
  .m_axi_rid      ( slave_slice_r_id         ),
  .m_axi_rdata    ( slave_slice[3].r_data    ),
  .m_axi_rresp    ( slave_slice[3].r_resp    ),
  .m_axi_rlast    ( slave_slice[3].r_last    ),
  .m_axi_rvalid   ( slave_slice[3].r_valid   ),
  .m_axi_rready   ( slave_slice[3].r_ready   ),
  // from size converter
  .s_axi_aclk     ( pcie_axi_clk             ),
  .s_axi_aresetn  ( ndmreset_n               ),
  .s_axi_awid     ( '0                       ),
  .s_axi_awaddr   ( pcie_dwidth_axi_awaddr   ),
  .s_axi_awlen    ( pcie_dwidth_axi_awlen    ),
  .s_axi_awsize   ( pcie_dwidth_axi_awsize   ),
  .s_axi_awburst  ( pcie_dwidth_axi_awburst  ),
  .s_axi_awlock   ( pcie_dwidth_axi_awlock   ),
  .s_axi_awcache  ( pcie_dwidth_axi_awcache  ),
  .s_axi_awprot   ( pcie_dwidth_axi_awprot   ),
  .s_axi_awregion ( pcie_dwidth_axi_awregion ),
  .s_axi_awqos    ( pcie_dwidth_axi_awqos    ),
  .s_axi_awvalid  ( pcie_dwidth_axi_awvalid  ),
  .s_axi_awready  ( pcie_dwidth_axi_awready  ),
  .s_axi_wdata    ( pcie_dwidth_axi_wdata    ),
  .s_axi_wstrb    ( pcie_dwidth_axi_wstrb    ),
  .s_axi_wlast    ( pcie_dwidth_axi_wlast    ),
  .s_axi_wvalid   ( pcie_dwidth_axi_wvalid   ),
  .s_axi_wready   ( pcie_dwidth_axi_wready   ),
  .s_axi_bid      (                          ),
  .s_axi_bresp    ( pcie_dwidth_axi_bresp    ),
  .s_axi_bvalid   ( pcie_dwidth_axi_bvalid   ),
  .s_axi_bready   ( pcie_dwidth_axi_bready   ),
  .s_axi_arid     ( '0                       ),
  .s_axi_araddr   ( pcie_dwidth_axi_araddr   ),
  .s_axi_arlen    ( pcie_dwidth_axi_arlen    ),
  .s_axi_arsize   ( pcie_dwidth_axi_arsize   ),
  .s_axi_arburst  ( pcie_dwidth_axi_arburst  ),
  .s_axi_arlock   ( pcie_dwidth_axi_arlock   ),
  .s_axi_arcache  ( pcie_dwidth_axi_arcache  ),
  .s_axi_arprot   ( pcie_dwidth_axi_arprot   ),
  .s_axi_arregion ( pcie_dwidth_axi_arregion ),
  .s_axi_arqos    ( pcie_dwidth_axi_arqos    ),
  .s_axi_arvalid  ( pcie_dwidth_axi_arvalid  ),
  .s_axi_arready  ( pcie_dwidth_axi_arready  ),
  .s_axi_rid      (                          ),
  .s_axi_rdata    ( pcie_dwidth_axi_rdata    ),
  .s_axi_rresp    ( pcie_dwidth_axi_rresp    ),
  .s_axi_rlast    ( pcie_dwidth_axi_rlast    ),
  .s_axi_rvalid   ( pcie_dwidth_axi_rvalid   ),
  .s_axi_rready   ( pcie_dwidth_axi_rready   )
);
`endif

endmodule
