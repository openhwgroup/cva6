// Copyright 2021 OpenHW Group
// Copyright 2021 Silicon Labs, Inc.
//
// Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     https://solderpad.org/licenses/
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


`include "uvma_isa_if.sv"


package uvma_isa_pkg;

  import uvm_pkg::*;
  import uvml_trn_pkg::*;

  `include "uvma_isa_cntxt.sv"
  `include "uvma_isa_mon_trn.sv"
  `include "uvma_isa_cov_model.sv"
  `include "uvma_isa_mon.sv"
  `include "uvma_isa_agent.sv"

endpackage : uvma_isa_pkg
