// COPYRIGHT HEADER


`ifndef __UVMA_RESET_IF_CHK_SV__
`define __UVMA_RESET_IF_CHK_SV__


/**
 * Encapsulates assertions targeting uvma_reset_if.
 */
module uvma_reset_if_chk(
   uvma_reset_if  reset_if
);
   
   `pragma protect begin
   
   // TODO Add assertions to uvma_reset_if_chk
   
   `pragma protect end
   
endmodule : uvma_reset_if_chk


`endif // __UVMA_RESET_IF_CHK_SV__
