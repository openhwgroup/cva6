/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 141;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000064,
        64'h65646E65_7478652D,
        64'h73747075_72726574,
        64'h6E690073_65676E61,
        64'h7200656C_646E6168,
        64'h70007265_6C6C6F72,
        64'h746E6F63_2D747075,
        64'h72726574_6E690073,
        64'h6C6C6563_2D747075,
        64'h72726574_6E692300,
        64'h79636E65_75716572,
        64'h662D6B63_6F6C6300,
        64'h65707974_2D756D6D,
        64'h00617369_2C766373,
        64'h69720073_75746174,
        64'h73006765_72006570,
        64'h79745F65_63697665,
        64'h64007963_6E657571,
        64'h6572662D_65736162,
        64'h656D6974_006C6564,
        64'h6F6D0065_6C626974,
        64'h61706D6F_6300736C,
        64'h6C65632D_657A6973,
        64'h2300736C_6C65632D,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_00000030,
        64'h66697468_2C626375,
        64'h1B000000_0A000000,
        64'h03000000_00000000,
        64'h66697468_01000000,
        64'h02000000_02000000,
        64'h00000C00_00000000,
        64'h00000002_00000000,
        64'h4B000000_10000000,
        64'h03000000_07000000,
        64'h01000000_03000000,
        64'h01000000_AE000000,
        64'h10000000_03000000,
        64'h00000000_30746E69,
        64'h6C632C76_63736972,
        64'h1B000000_0D000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6E696C63_01000000,
        64'hA7000000_00000000,
        64'h03000000_00007375,
        64'h622D656C_706D6973,
        64'h00636F73_2D657261,
        64'h622D656E_61697261,
        64'h2C687465_1B000000,
        64'h1F000000_03000000,
        64'h02000000_0F000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636F73_01000000,
        64'h02000000_00000001,
        64'h00000000_00000080,
        64'h00000000_4B000000,
        64'h10000000_03000000,
        64'h00007972_6F6D656D,
        64'h3F000000_07000000,
        64'h03000000_00303030,
        64'h30303030_38407972,
        64'h6F6D656D_01000000,
        64'h02000000_02000000,
        64'h02000000_01000000,
        64'h9F000000_04000000,
        64'h03000000_00006374,
        64'h6E692D75_70632C76,
        64'h63736972_1B000000,
        64'h0F000000_03000000,
        64'h8A000000_00000000,
        64'h03000000_01000000,
        64'h79000000_04000000,
        64'h03000000_00000000,
        64'h72656C6C_6F72746E,
        64'h6F632D74_70757272,
        64'h65746E69_01000000,
        64'h00CA9A3B_69000000,
        64'h04000000_03000000,
        64'h00003933_76732C76,
        64'h63736972_60000000,
        64'h0B000000_03000000,
        64'h00636D69_34367672,
        64'h56000000_08000000,
        64'h03000000_00000076,
        64'h63736972_1B000000,
        64'h06000000_03000000,
        64'h00000000_79616B6F,
        64'h4F000000_05000000,
        64'h03000000_00000000,
        64'h4B000000_04000000,
        64'h03000000_00757063,
        64'h3F000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h80969800_2C000000,
        64'h04000000_03000000,
        64'h00000000_0F000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_00657261,
        64'h622D656E_61697261,
        64'h2C687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2D657261,
        64'h622D656E_61697261,
        64'h2C687465_1B000000,
        64'h14000000_03000000,
        64'h02000000_0F000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hE8020000_C2000000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h20030000_38000000,
        64'hE2030000_EDFE0DD0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_0000BFF5,
        64'h10500073_03C58593,
        64'h00000597_F1402573,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00008402_07458593,
        64'h00000597_F1402573,
        64'h01F41413_0010041B
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into 
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q<RomSize) ? mem[addr_q] : '0;
endmodule
