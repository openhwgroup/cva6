///////////////////////////////////////////////////////////////////////////////
//
// Copyright 2021 OpenHW Group
// Copyright 2021 Thales DIS Design Services SAS
//
// Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//    https://solderpad.org/licenses/
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.0
//
///////////////////////////////////////////////////////////////////////////////
//
// CVA6 "core_only" testbench wrapper.
//
///////////////////////////////////////////////////////////////////////////////

`define MAIN_MEM(P) uvmt_cva6_tb.cva6_dut_wrap.cva6_tb_wrapper_i.i_sram.gen_cut[0].gen_mem.i_tc_sram_wrapper.i_tc_sram.init_val[(``P``)]
`define USER_MEM(P) uvmt_cva6_tb.cva6_dut_wrap.cva6_tb_wrapper_i.i_sram.gen_cut[0].gen_mem.gen_mem_user.i_tc_sram_wrapper_user.i_tc_sram.init_val[(``P``)]

import uvm_pkg::*;

`include "uvm_macros.svh"

import "DPI-C" function read_elf(input string filename);
import "DPI-C" function byte get_section(output longint address, output longint len);
import "DPI-C" context function void read_section(input longint address, inout byte buffer[]);

module cva6_tb_wrapper #(
  parameter int unsigned AXI_USER_WIDTH    = 1,
  parameter int unsigned AXI_USER_EN       = 0,
  parameter int unsigned AXI_ADDRESS_WIDTH = 64,
  parameter int unsigned AXI_DATA_WIDTH    = 64,
  parameter int unsigned NUM_WORDS         = 2**25
) (
  input  logic                         clk_i,
  input  logic                         rst_ni,
  output wire                          tb_exit_o,
  output ariane_rvfi_pkg::rvfi_port_t  rvfi_o,
  input  cvxif_pkg::cvxif_resp_t       cvxif_resp,
  output cvxif_pkg::cvxif_req_t        cvxif_req,
  uvma_axi_intf                        axi_slave
);

  ariane_axi::req_t    axi_ariane_req;
  ariane_axi::resp_t   axi_ariane_resp;

  static uvm_cmdline_processor uvcl = uvm_cmdline_processor::get_inst();
  string binary = "";

  ariane_rvfi_pkg::rvfi_port_t  rvfi;
  assign rvfi_o = rvfi;

  cva6 #(
    .ArianeCfg  ( ariane_soc::ArianeSocCfg )
  ) i_cva6 (
    .clk_i                ( clk_i                     ),
    .rst_ni               ( rst_ni                    ),
    .boot_addr_i          ( 64'h0000_0000_8000_0000   ), //ariane_soc::ROMBase
    .hart_id_i            ( 64'h0000_0000_0000_0000   ),
    .irq_i                ( 2'b00 /*irqs*/            ),
    .ipi_i                ( 1'b0  /*ipi*/             ),
    .time_irq_i           ( 1'b0  /*timer_irq*/       ),
    .debug_req_i          ( 1'b0                      ),
    .rvfi_o               ( rvfi                      ),
    .cvxif_req_o          ( cvxif_req                 ),
    .cvxif_resp_i         ( cvxif_resp                ),
    .axi_req_o            ( axi_ariane_req            ),
    .axi_resp_i           ( axi_ariane_resp           )
  );

  //----------------------------------------------------------------------------
  // RVFI
  //----------------------------------------------------------------------------

  rvfi_tracer  #(
    .HART_ID(8'h0),
    .DEBUG_START(0),
    .DEBUG_STOP(0),
    .NR_COMMIT_PORTS(ariane_pkg::NR_COMMIT_PORTS)
  ) rvfi_tracer_i (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .rvfi_i(rvfi)
  ) ;

  //----------------------------------------------------------------------------
  // Memory
  //----------------------------------------------------------------------------

  logic                         req;
  logic                         we;
  logic [AXI_ADDRESS_WIDTH-1:0] addr;
  logic [AXI_DATA_WIDTH/8-1:0]  be;
  logic [AXI_DATA_WIDTH-1:0]    wdata;
  logic [AXI_USER_WIDTH-1:0]    wuser;
  logic [AXI_DATA_WIDTH-1:0]    rdata;
  logic [AXI_USER_WIDTH-1:0]    ruser;

  AXI_BUS #(
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH        ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH           ),
    .AXI_ID_WIDTH   ( ariane_soc::IdWidthSlave ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH           )
  ) cva6_axi_bus();

  axi_master_connect #(
  ) i_axi_master_connect_cva6_to_mem (
    .axi_req_i  (axi_ariane_req),
    .axi_resp_o (axi_ariane_resp),
    .master     (cva6_axi_bus)
  );

  axi2mem #(
    .AXI_ID_WIDTH   ( ariane_soc::IdWidthSlave ),
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH        ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH           ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH           )
  ) i_cva6_axi2mem (
    .clk_i  ( clk_i       ),
    .rst_ni ( rst_ni      ),
    .slave  ( cva6_axi_bus ),
    .req_o  ( req          ),
    .we_o   ( we           ),
    .addr_o ( addr         ),
    .be_o   ( be           ),
    .user_o ( wuser        ),
    .data_o ( wdata        ),
    .user_i ( ruser        ),
    .data_i ( rdata        )
  );

  sram #(
    .USER_WIDTH ( AXI_USER_WIDTH ),
    .DATA_WIDTH ( AXI_DATA_WIDTH ),
    .USER_EN    ( AXI_USER_EN    ),
    .SIM_INIT   ( "zeros"        ),
    .NUM_WORDS  ( NUM_WORDS      )
  ) i_sram (
    .clk_i      ( clk_i                                                                       ),
    .rst_ni     ( rst_ni                                                                      ),
    .req_i      ( req                                                                         ),
    .we_i       ( we                                                                          ),
    .addr_i     ( addr[$clog2(NUM_WORDS)-1+$clog2(AXI_DATA_WIDTH/8):$clog2(AXI_DATA_WIDTH/8)] ),
    .wuser_i    ( wuser                                                                       ),
    .wdata_i    ( wdata                                                                       ),
    .be_i       ( be                                                                          ),
    .ruser_o    ( ruser                                                                       ),
    .rdata_o    ( rdata                                                                       )
  );

   // AW Channel
   assign axi_slave.aw_valid  = cva6_axi_bus.aw_valid;
   assign axi_slave.aw_ready  = cva6_axi_bus.aw_ready;
   assign axi_slave.aw_id     = cva6_axi_bus.aw_id;
   assign axi_slave.aw_addr   = cva6_axi_bus.aw_addr;
   assign axi_slave.aw_len    = cva6_axi_bus.aw_len;
   assign axi_slave.aw_size   = cva6_axi_bus.aw_size;
   assign axi_slave.aw_burst  = cva6_axi_bus.aw_burst;
   assign axi_slave.aw_lock   = cva6_axi_bus.aw_lock;
   assign axi_slave.aw_cache  = cva6_axi_bus.aw_cache;
   assign axi_slave.aw_prot   = cva6_axi_bus.aw_prot;
   assign axi_slave.aw_qos    = cva6_axi_bus.aw_qos;
   assign axi_slave.aw_region = cva6_axi_bus.aw_region;
   assign axi_slave.aw_user   = cva6_axi_bus.aw_user;
   assign axi_slave.aw_atop   = cva6_axi_bus.aw_atop;
   // W Channel
   assign axi_slave.w_valid = cva6_axi_bus.w_valid;
   assign axi_slave.w_ready = cva6_axi_bus.w_ready;
   assign axi_slave.w_data  = cva6_axi_bus.w_data;
   assign axi_slave.w_strb  = cva6_axi_bus.w_strb;
   assign axi_slave.w_last  = cva6_axi_bus.w_last;
   assign axi_slave.w_user  = cva6_axi_bus.w_user;
   // B Channel
   assign axi_slave.b_valid = cva6_axi_bus.b_valid;
   assign axi_slave.b_ready = cva6_axi_bus.b_ready;
   assign axi_slave.b_id    = cva6_axi_bus.b_id;
   assign axi_slave.b_resp  = cva6_axi_bus.b_resp;
   assign axi_slave.b_user  = cva6_axi_bus.b_user;
   // AR Channel
   assign axi_slave.ar_valid  = cva6_axi_bus.ar_valid;
   assign axi_slave.ar_ready  = cva6_axi_bus.ar_ready;
   assign axi_slave.ar_id     = cva6_axi_bus.ar_id;
   assign axi_slave.ar_addr   = cva6_axi_bus.ar_addr;
   assign axi_slave.ar_len    = cva6_axi_bus.ar_len;
   assign axi_slave.ar_size   = cva6_axi_bus.ar_size;
   assign axi_slave.ar_burst  = cva6_axi_bus.ar_burst;
   assign axi_slave.ar_lock   = cva6_axi_bus.ar_lock;
   assign axi_slave.ar_cache  = cva6_axi_bus.ar_cache;
   assign axi_slave.ar_prot   = cva6_axi_bus.ar_prot;
   assign axi_slave.ar_qos    = cva6_axi_bus.ar_qos;
   assign axi_slave.ar_region = cva6_axi_bus.ar_region;
   assign axi_slave.ar_user   = cva6_axi_bus.ar_user;
   // R Channel
   assign axi_slave.r_valid = cva6_axi_bus.r_valid;
   assign axi_slave.r_ready = cva6_axi_bus.r_ready;
   assign axi_slave.r_id    = cva6_axi_bus.r_id;
   assign axi_slave.r_data  = cva6_axi_bus.r_data;
   assign axi_slave.r_resp  = cva6_axi_bus.r_resp;
   assign axi_slave.r_last  = cva6_axi_bus.r_last;
   assign axi_slave.r_user  = cva6_axi_bus.r_user;
    initial begin
        automatic logic [7:0][7:0] mem_row;
        longint address;
        longint len;
        byte buffer[];
        void'(uvcl.get_arg_value("+PRELOAD=", binary));

        if (binary != "") begin

            void'(read_elf(binary));

            wait(clk_i);

            // while there are more sections to process
            while (get_section(address, len)) begin
                automatic int num_words0 = (len+7)/8;
                `uvm_info( "Core Test", $sformatf("Loading Address: %x, Length: %x", address, len), UVM_LOW)
                buffer = new [num_words0*8];
                void'(read_section(address, buffer));
                // preload memories
                // 64-bit
                for (int i = 0; i < num_words0; i++) begin
                    mem_row = '0;
                    for (int j = 0; j < 8; j++) begin
                        mem_row[j] = buffer[i*8 + j];
                    end
                    `MAIN_MEM((address[23:0] >> 3) + i) = mem_row;
                end
            end
        end
    end

endmodule
