// COPYRIGHT HEADER


`ifndef __UVML_LOGS_TDEFS_SV__
`define __UVML_LOGS_TDEFS_SV__





`endif // __UVML_LOGS_TDEFS_SV__
