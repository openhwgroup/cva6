package alu_sequence_pkg;


import fu_if_agent_pkg::*;
import uvm_pkg::*;
import ariane_pkg::*;

`include "uvm_macros.svh"
`include "fibonacci_sequence.svh"
`include "reset_sequence.svh"
`include "basic_sequence.svh"
`include "add_sequence.svh"
`include "addw_sequence.svh"
`include "subw_sequence.svh"
`include "sub_sequence.svh"
`include "xor_sequence.svh"
`include "or_sequence.svh"
`include "and_sequence.svh"

endpackage
