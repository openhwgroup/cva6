/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 1024;

    const logic [RomSize-1:0][31:0] mem_H = {
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h0a0d2165,
        32'h00000000,
        32'h616d6920,
        32'h20676e69,
        32'h00000000,
        32'h3a656d61,
        32'h00093a73,
        32'h69727474,
        32'h00000009,
        32'h20747361,
        32'h0000093a,
        32'h74737269,
        32'h00000000,
        32'h09202020,
        32'h69756720,
        32'h69747261,
        32'h00000000,
        32'h093a6469,
        32'h70797420,
        32'h69747261,
        32'h00000000,
        32'h6e65206e,
        32'h74726170,
        32'h00000009,
        32'h65697274,
        32'h6f697469,
        32'h20657a69,
        32'h00000009,
        32'h72746e65,
        32'h74697472,
        32'h65626d75,
        32'h00000009,
        32'h61626c20,
        32'h746e6520,
        32'h69747261,
        32'h00093a61,
        32'h756b6361,
        32'h00000000,
        32'h093a6162,
        32'h65727275,
        32'h00000009,
        32'h72657365,
        32'h00093a72,
        32'h685f6372,
        32'h00000000,
        32'h3a657a69,
        32'h00000009,
        32'h73697665,
        32'h0000093a,
        32'h616e6769,
        32'h00000000,
        32'h64616568,
        32'h6174206e,
        32'h74726170,
        32'h0000203a,
        32'h76206e72,
        32'h2079706f,
        32'h00000000,
        32'h0d216465,
        32'h20647261,
        32'h00000000,
        32'h0d216465,
        32'h6974696e,
        32'h00000000,
        32'h69746978,
        32'h2e647320,
        32'h61697469,
        32'h6f6e2064,
        32'h00000000,
        32'h00000000,
        32'h0d6b636f,
        32'h53206461,
        32'h6f6e2064,
        32'h0000000a,
        32'h2e445320,
        32'h696c6169,
        32'h00000031,
        32'h00000035,
        32'h00000000,
        32'h00000020,
        32'h6e6f7073,
        32'h00000000,
        32'h616d6d6f,
        32'h00000000,
        32'h74706d65,
        32'h206f6669,
        32'h00000000,
        32'h2164657a,
        32'h74696e69,
        32'h00000000,
        32'h203a7375,
        32'h00000000,
        32'h49505320,
        32'h00000a0d,
        32'h6f57206f,
        32'h00000000,
        32'h2d746c75,
        32'h2d697274,
        32'h7800746c,
        32'h642d6972,
        32'h6c78006c,
        32'h73692c78,
        32'h746e6573,
        32'h74707572,
        32'h692c786e,
        32'h74646977,
        32'h70672c78,
        32'h68746469,
        32'h70672c78,
        32'h322d746c,
        32'h642d7475,
        32'h6e6c7800,
        32'h6665642d,
        32'h2c786e6c,
        32'h73747570,
        32'h6c612c78,
        32'h73747570,
        32'h6c612c78,
        32'h72656c6c,
        32'h6f632d6f,
        32'h736c6c65,
        32'h70672300,
        32'h6464612d,
        32'h6c61636f,
        32'h2d656c62,
        32'h00736567,
        32'h65676174,
        32'h79636e65,
        32'h662d7861,
        32'h73006f69,
        32'h6b63732c,
        32'h00737469,
        32'h66736e61,
        32'h756e2c78,
        32'h73746962,
        32'h6d756e2c,
        32'h00747369,
        32'h6669662c,
        32'h00796c69,
        32'h786e6c78,
        32'h69772d6f,
        32'h72007466,
        32'h67657200,
        32'h72726574,
        32'h6e657261,
        32'h75727265,
        32'h64656570,
        32'h65727275,
        32'h646e2c76,
        32'h00797469,
        32'h702d7861,
        32'h73697200,
        32'h6e2d6765,
        32'h646e6574,
        32'h74707572,
        32'h69007365,
        32'h00646564,
        32'h75732d65,
        32'h2d6e6961,
        32'h72656767,
        32'h746c7561,
        32'h78756e69,
        32'h69706700,
        32'h61687000,
        32'h6f72746e,
        32'h70757272,
        32'h00736c6c,
        32'h70757272,
        32'h23007469,
        32'h626c7400,
        32'h2d756d6d,
        32'h2c766373,
        32'h75746174,
        32'h72006570,
        32'h63697665,
        32'h6e657571,
        32'h6b636f6c,
        32'h6e657571,
        32'h65736162,
        32'h00687461,
        32'h6f647473,
        32'h6f6d0065,
        32'h61706d6f,
        32'h6c65632d,
        32'h2300736c,
        32'h73736572,
        32'h09000000,
        32'h02000000,
        32'h01000000,
        32'h04000000,
        32'hffffffff,
        32'h04000000,
        32'hffffffff,
        32'h04000000,
        32'h01000000,
        32'h04000000,
        32'h00000000,
        32'h04000000,
        32'h08000000,
        32'h04000000,
        32'h08000000,
        32'h04000000,
        32'h00000000,
        32'h04000000,
        32'h00000000,
        32'h04000000,
        32'h00000000,
        32'h04000000,
        32'h00000000,
        32'h04000000,
        32'h00000100,
        32'h00000040,
        32'h67000000,
        32'h03000000,
        32'h00000000,
        32'h00000000,
        32'h2e312d6f,
        32'h7370782c,
        32'h1b000000,
        32'h03000000,
        32'h05020000,
        32'h03000000,
        32'h30303030,
        32'h6f697067,
        32'h02000000,
        32'h00000000,
        32'h00000000,
        32'h10000000,
        32'h00007fe3,
        32'hf3010000,
        32'h03000000,
        32'h03000000,
        32'h08000000,
        32'h03000000,
        32'h04000000,
        32'h006b726f,
        32'h5b000000,
        32'h03000000,
        32'h2d637369,
        32'h1b000000,
        32'h03000000,
        32'h30303030,
        32'h40687465,
        32'h72776f6c,
        32'h02000000,
        32'he8010000,
        32'h03000000,
        32'he40c0000,
        32'h08000000,
        32'h20bcbe00,
        32'h04000000,
        32'h00000000,
        32'h04000000,
        32'h00000000,
        32'h2d697073,
        32'h1b000000,
        32'h03000000,
        32'h40636d6d,
        32'h04000000,
        32'h04000000,
        32'h08000000,
        32'h04000000,
        32'h01000000,
        32'h04000000,
        32'h01000000,
        32'h04000000,
        32'h00377865,
        32'h74010000,
        32'h03000000,
        32'h00000000,
        32'h00000000,
        32'h10000000,
        32'h02000000,
        32'h52010000,
        32'h03000000,
        32'h41010000,
        32'h03000000,
        32'h0f000000,
        32'h03000000,
        32'h00000000,
        32'h03000000,
        32'h302e322d,
        32'h7370782c,
        32'h00622e30,
        32'h6970732d,
        32'h786e6c78,
        32'h28000000,
        32'h00000000,
        32'h30303032,
        32'h2d737078,
        32'h02000000,
        32'h67010000,
        32'h03000000,
        32'h5d010000,
        32'h03000000,
        32'h52010000,
        32'h03000000,
        32'h41010000,
        32'h03000000,
        32'h33010000,
        32'h03000000,
        32'h4b000000,
        32'h03000000,
        32'h00000000,
        32'h00000000,
        32'h10000000,
        32'h00303537,
        32'h1b000000,
        32'h03000000,
        32'h30303030,
        32'h74726175,
        32'h02000000,
        32'h746e6f63,
        32'h08000000,
        32'h00100000,
        32'h00000000,
        32'h67000000,
        32'h03000000,
        32'h02000000,
        32'h08000000,
        32'h00333130,
        32'h65642c76,
        32'h1b000000,
        32'h03000000,
        32'h72656c6c,
        32'h6f632d67,
        32'h01000000,
        32'h03000000,
        32'h04000000,
        32'h03000000,
        32'h04000000,
        32'h07000000,
        32'h04000000,
        32'h00000004,
        32'h0000000c,
        32'h67000000,
        32'h03000000,
        32'h02000000,
        32'h02000000,
        32'h10000000,
        32'ha0000000,
        32'h03000000,
        32'h6c702c76,
        32'h1b000000,
        32'h03000000,
        32'h8f000000,
        32'h03000000,
        32'h00000000,
        32'h03000000,
        32'h30303030,
        32'h72656c6c,
        32'h6f632d74,
        32'h65746e69,
        32'h02000000,
        32'h746e6f63,
        32'h08000000,
        32'h00000c00,
        32'h00000002,
        32'h67000000,
        32'h03000000,
        32'h02000000,
        32'h02000000,
        32'h10000000,
        32'h00000000,
        32'h6c632c76,
        32'h1b000000,
        32'h03000000,
        32'h30303030,
        32'h6e696c63,
        32'hf0000000,
        32'h03000000,
        32'h622d656c,
        32'h00636f73,
        32'h622d656e,
        32'h2c687465,
        32'h1f000000,
        32'h02000000,
        32'h04000000,
        32'h02000000,
        32'h04000000,
        32'h00636f73,
        32'h02000000,
        32'hd9000000,
        32'h03000000,
        32'h61656274,
        32'hc3000000,
        32'h03000000,
        32'h01000000,
        32'hbd000000,
        32'h03000000,
        32'h656c2d74,
        32'h72616568,
        32'h00000073,
        32'h6f697067,
        32'h0a000000,
        32'h00000000,
        32'h01000000,
        32'h00000040,
        32'h00000080,
        32'h67000000,
        32'h03000000,
        32'h6f6d656d,
        32'h07000000,
        32'h00303030,
        32'h38407972,
        32'h01000000,
        32'h02000000,
        32'h02000000,
        32'h04000000,
        32'h00006374,
        32'h70632c76,
        32'h1b000000,
        32'h03000000,
        32'h00000000,
        32'h01000000,
        32'h04000000,
        32'h00000000,
        32'h6f72746e,
        32'h70757272,
        32'h01000000,
        32'h00000000,
        32'h00003933,
        32'h63736972,
        32'h0b000000,
        32'h00006364,
        32'h34367672,
        32'h0b000000,
        32'h00000076,
        32'h00656e61,
        32'h2c687465,
        32'h12000000,
        32'h00000000,
        32'h6b000000,
        32'h03000000,
        32'h67000000,
        32'h03000000,
        32'h5b000000,
        32'h03000000,
        32'h4b000000,
        32'h03000000,
        32'h40757063,
        32'hc0e1e400,
        32'h04000000,
        32'h00000000,
        32'h04000000,
        32'h01000000,
        32'h04000000,
        32'h00000000,
        32'h01000000,
        32'h00000030,
        32'h313a3030,
        32'h30314074,
        32'h636f732f,
        32'h1a000000,
        32'h00006e65,
        32'h01000000,
        32'h622d656e,
        32'h2c687465,
        32'h10000000,
        32'h00766564,
        32'h622d656e,
        32'h2c687465,
        32'h14000000,
        32'h02000000,
        32'h04000000,
        32'h02000000,
        32'h04000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'hd0080000,
        32'h00000000,
        32'h11000000,
        32'h08090000,
        32'hda0b0000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h46454443,
        32'h37363534,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h13058593,
        32'h01f41413,
        32'he911d05f,
        32'h65a14505,
        32'hd3050513,
        32'he84ff0ef,
        32'h05132005,
        32'h02faf537,
        32'hee0ff0ef,
        32'h00001517,
        32'h05130000,
        32'hf0ef8526,
        32'hea050513,
        32'hf08ff0ef,
        32'h00001517,
        32'h05130000,
        32'hf0ef8526,
        32'hec850513,
        32'hf30ff0ef,
        32'h00001517,
        32'hc3dff0ef,
        32'h020b2583,
        32'h09850513,
        32'hf3849de3,
        32'h080a0993,
        32'h2485e1a5,
        32'h1517ff3a,
        32'hf0ef0a05,
        32'hf80ff0ef,
        32'h00001517,
        32'h01093503,
        32'h0c050513,
        32'h823ff0ef,
        32'hfa8ff0ef,
        32'h00001517,
        32'hfb898a13,
        32'hfc0ff0ef,
        32'h00001517,
        32'h895ff0ef,
        32'h4503f909,
        32'hf0ef0ca5,
        32'h1517ff9a,
        32'hf0ef0a05,
        32'h014d07b3,
        32'hf0eff809,
        32'h05130000,
        32'hf0ef0ff4,
        32'hf0ef0ca5,
        32'h15174c11,
        32'h1b630201,
        32'h099384aa,
        32'hf0ef850a,
        32'h04892583,
        32'hef850513,
        32'h893ff0ef,
        32'hf0ef0ea5,
        32'h15178a5f,
        32'h869ff0ef,
        32'h00001517,
        32'h652687bf,
        32'h05130000,
        32'hf0ef7502,
        32'h0d050513,
        32'h91bff0ef,
        32'hf0ef0ca5,
        32'h15178edf,
        32'h8b1ff0ef,
        32'h00001517,
        32'h45428c3f,
        32'h05130000,
        32'hf0ef4532,
        32'h0d050513,
        32'h923ff0ef,
        32'hf0ef0d25,
        32'h1517975f,
        32'h8f9ff0ef,
        32'h00001517,
        32'h0c050513,
        32'hbf5154f9,
        32'hfc850513,
        32'h9a3ff0ef,
        32'hf0ef0ca5,
        32'h1517933f,
        32'h05130000,
        32'h84aa890a,
        32'h850a4585,
        32'h951ff0ef,
        32'h00001517,
        32'h6d026ca2,
        32'h7b027aa2,
        32'h690664a6,
        32'h60e6fa04,
        32'h981ff0ef,
        32'h00001517,
        32'hf0ef8bae,
        32'he06ae466,
        32'hf852fc4e,
        32'hec86ec5e,
        32'h711db765,
        32'h61696baa,
        32'h7a0a79aa,
        32'h640e60ae,
        32'h9d1ff0ef,
        32'h00001517,
        32'hc61ff0ef,
        32'hc69ff0ef,
        32'hc71ff0ef,
        32'hc79ff0ef,
        32'hf0efc8bf,
        32'h45814605,
        32'h46e32004,
        32'ha19ff0ef,
        32'h00001517,
        32'he7b30689,
        32'h29011442,
        32'hf0ef9041,
        32'h0085151b,
        32'hfc941ae3,
        32'hff7a17e3,
        32'hf0ef0a05,
        32'hc5830144,
        32'h0b934a01,
        32'h850a0400,
        32'h4901ff55,
        32'hf0efe004,
        32'h0b130fe0,
        32'h20048493,
        32'h454985a2,
        32'h00166613,
        32'hf4dff0ef,
        32'hf55ff0ef,
        32'h0084559b,
        32'h0ff5f593,
        32'hf6dff0ef,
        32'h559bfee7,
        32'h00c68023,
        32'h08000713,
        32'h0209d993,
        32'he55ee95a,
        32'hf94ae586,
        32'h02061993,
        32'h80829141,
        32'h8ff90057,
        32'h67090107,
        32'h179b4105,
        32'h151b8d2d,
        32'h8da9893d,
        32'h8da99141,
        32'h05220085,
        32'h07f57513,
        32'h15938d2d,
        32'hd51b0075,
        32'h80820141,
        32'h60a257f5,
        32'hf89ff0ef,
        32'hefbff0ef,
        32'heb7ff0ef,
        32'hf0ef347d,
        32'hf0ef29a5,
        32'h1517c89f,
        32'he4061141,
        32'h00153513,
        32'h60e20004,
        32'h0ce3e3bf,
        32'hf0ef2c25,
        32'h151785aa,
        32'hf0ef0290,
        32'h05b70770,
        32'hf0ef4485,
        32'he4261101,
        32'h00153513,
        32'h60a20004,
        32'hf0ef2fc5,
        32'h00001517,
        32'h842ae9bf,
        32'he4060370,
        32'h06500613,
        32'h61056902,
        32'h60e20015,
        32'h05130004,
        32'h986388bd,
        32'h45014785,
        32'hed1ff0ef,
        32'hf0ef84aa,
        32'hee1ff0ef,
        32'h892aef3f,
        32'he426e822,
        32'h1aa00593,
        32'h1101bfcd,
        32'h61056902,
        32'h60e24505,
        32'h458538a5,
        32'h1517fe99,
        32'hf29ff0ef,
        32'hf39ff0ef,
        32'h09500613,
        32'h0413e04a,
        32'h6409e822,
        32'hf06f6105,
        32'h00001517,
        32'hda5ff0ef,
        32'hce9ff0ef,
        32'h00001517,
        32'h8522cfbf,
        32'hec063d25,
        32'h1517842a,
        32'h80826145,
        32'h70a2f47d,
        32'hd4634187,
        32'h179bfabf,
        32'hf0ef8532,
        32'h6622ec1f,
        32'h7513ec9f,
        32'h75130084,
        32'hf0ef0ff5,
        32'h551bee1f,
        32'h551bee9f,
        32'he513febf,
        32'h842eec26,
        32'hf4067179,
        32'h0ff00513,
        32'hb7d900d7,
        32'h00f60733,
        32'hff698b05,
        32'hd6b80785,
        32'h00f50733,
        32'hd3b84719,
        32'h200007b7,
        32'h0007869b,
        32'h20000537,
        32'h537c2000,
        32'h200007b7,
        32'hfff537fd,
        32'h079304b7,
        32'h871b4781,
        32'hdbb85779,
        32'h06b7ee63,
        32'h80826105,
        32'h4719dbb8,
        32'h0ff47513,
        32'h07b7e23f,
        32'h05130000,
        32'hf0ef9101,
        32'he39ff0ef,
        32'h00001517,
        32'h240153fc,
        32'h8b050647,
        32'hd3b81060,
        32'h07b7fff5,
        32'h06400793,
        32'h5779e426,
        32'h200007b7,
        32'hf06f6105,
        32'h00001517,
        32'h6442d03c,
        32'hf0ef54a5,
        32'h1517f25f,
        32'h02049513,
        32'hf0ef5425,
        32'h15175064,
        32'h0793ec3f,
        32'h05130000,
        32'hf0ef9101,
        32'h2481edbf,
        32'h05130000,
        32'hd03c1040,
        32'h0437fff5,
        32'h47a9c3b8,
        32'h07b7f03f,
        32'he822ec06,
        32'h11010000,
        32'h25014108,
        32'h80826105,
        32'hf0ef0091,
        32'hf0ef0081,
        32'hf0efec06,
        32'h80826145,
        32'h740270a2,
        32'hef9ff0ef,
        32'hf01ff0ef,
        32'h4503f81f,
        32'h7513002c,
        32'h54e10380,
        32'hf406e84a,
        32'h71798082,
        32'h64e27402,
        32'h10e3f3bf,
        32'h4503f43f,
        32'h00814503,
        32'h0ff57513,
        32'h553b54e1,
        32'hf406e84a,
        32'h71798082,
        32'h0007c783,
        32'h97aa8111,
        32'h973e00f5,
        32'h87930000,
        32'h0405f93f,
        32'h01416402,
        32'h00044503,
        32'he0221141,
        32'h88230200,
        32'h8423fc70,
        32'h8623470d,
        32'h0ff57513,
        32'h0085551b,
        32'h00e78623,
        32'h00078223,
        32'h02b5553b,
        32'h808200a7,
        32'h0207f793,
        32'h10000737,
        32'h75130147,
        32'h07b78082,
        32'h808200b5,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00048067,
        32'h0010049b,
        32'h00001597,
        32'hff24c6e3,
        32'h02000937,
        32'hfe091ee3,
        32'h00092023,
        32'h00291913,
        32'h020004b7,
        32'h00897913,
        32'h10500073,
        32'h4009091b,
        32'h00448493,
        32'h00100913,
        32'h27f000ef,
        32'h0210011b,
        32'hf1402973,
        32'h30491073
    };

    const logic [RomSize-1:0][31:0] mem_L = {
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h6e6f6420,
        32'h00206567,
        32'h746f6f62,
        32'h79706f63,
        32'h00000009,
        32'h6e090a0d,
        32'h65747562,
        32'h61090a0d,
        32'h3a61626c,
        32'h6c090a0d,
        32'h61626c20,
        32'h66090a0d,
        32'h00000000,
        32'h20203a64,
        32'h6e6f6974,
        32'h70090a0d,
        32'h00000000,
        32'h75672065,
        32'h6e6f6974,
        32'h70090a0d,
        32'h20797274,
        32'h6f697469,
        32'h20747067,
        32'h20203a73,
        32'h6e65206e,
        32'h74726170,
        32'h73090a0d,
        32'h3a736569,
        32'h206e6f69,
        32'h61702072,
        32'h6e090a0d,
        32'h2020203a,
        32'h73656972,
        32'h6e6f6974,
        32'h70090a0d,
        32'h646c2070,
        32'h62090a0d,
        32'h00000000,
        32'h6c20746e,
        32'h63090a0d,
        32'h3a646576,
        32'h72090a0d,
        32'h65646165,
        32'h63090a0d,
        32'h00000909,
        32'h73090a0d,
        32'h3a6e6f69,
        32'h72090a0d,
        32'h65727574,
        32'h73090a0d,
        32'h003a7265,
        32'h20656c62,
        32'h6f697469,
        32'h20747067,
        32'h65756c61,
        32'h75746572,
        32'h63206473,
        32'h0000000a,
        32'h6c696166,
        32'h63204453,
        32'h0000000a,
        32'h7a696c61,
        32'h69206473,
        32'h0a0d676e,
        32'h65202e2e,
        32'h657a696c,
        32'h6e692074,
        32'h6c756f63,
        32'h0000002e,
        32'h0000000a,
        32'h6c622044,
        32'h65722074,
        32'h6c756f63,
        32'h0d202e2e,
        32'h676e697a,
        32'h74696e69,
        32'h34646d63,
        32'h35646d63,
        32'h30646d63,
        32'h3a206573,
        32'h65720920,
        32'h0020646e,
        32'h63204453,
        32'h203f3f79,
        32'h20746f6e,
        32'h66207872,
        32'h00000a0d,
        32'h696c6169,
        32'h20495053,
        32'h00007830,
        32'h74617473,
        32'h00000a0d,
        32'h74696e69,
        32'h21646c72,
        32'h6c6c6548,
        32'h00000032,
        32'h61666564,
        32'h2c786e6c,
        32'h75616665,
        32'h742c786e,
        32'h6175642d,
        32'h6e6c7800,
        32'h6572702d,
        32'h7265746e,
        32'h6c780068,
        32'h2d326f69,
        32'h6e6c7800,
        32'h772d6f69,
        32'h6e6c7800,
        32'h75616665,
        32'h6f642c78,
        32'h746c7561,
        32'h74756f64,
        32'h7800322d,
        32'h6e692d6c,
        32'h6e6c7800,
        32'h6e692d6c,
        32'h6e6c7800,
        32'h6f72746e,
        32'h69706700,
        32'h632d6f69,
        32'h73736572,
        32'h63616d2d,
        32'h6c007077,
        32'h61736964,
        32'h6e61722d,
        32'h6c6f7600,
        32'h75716572,
        32'h6d2d6970,
        32'h7461722d,
        32'h786e6c78,
        32'h622d7265,
        32'h72742d6d,
        32'h6e6c7800,
        32'h2d73732d,
        32'h786e6c78,
        32'h78652d6f,
        32'h786e6c78,
        32'h6d61662c,
        32'h00687464,
        32'h692d6765,
        32'h6968732d,
        32'h73747075,
        32'h6e690074,
        32'h702d7470,
        32'h746e6900,
        32'h732d746e,
        32'h63007665,
        32'h63736972,
        32'h726f6972,
        32'h6d2c7663,
        32'h73656d61,
        32'h72006465,
        32'h78652d73,
        32'h7265746e,
        32'h676e6172,
        32'h6e657073,
        32'h74617473,
        32'h74657200,
        32'h6972742d,
        32'h6665642c,
        32'h6c00736f,
        32'h656c646e,
        32'h72656c6c,
        32'h6f632d74,
        32'h65746e69,
        32'h65632d74,
        32'h65746e69,
        32'h6c70732d,
        32'h65707974,
        32'h00617369,
        32'h69720073,
        32'h73006765,
        32'h79745f65,
        32'h64007963,
        32'h6572662d,
        32'h63007963,
        32'h6572662d,
        32'h656d6974,
        32'h702d7475,
        32'h006c6564,
        32'h6c626974,
        32'h6300736c,
        32'h657a6973,
        32'h6c65632d,
        32'h64646123,
        32'h02000000,
        32'h02000000,
        32'hb5000000,
        32'h03000000,
        32'hbf020000,
        32'h03000000,
        32'hae020000,
        32'h03000000,
        32'ha1020000,
        32'h03000000,
        32'h8a020000,
        32'h03000000,
        32'h79020000,
        32'h03000000,
        32'h69020000,
        32'h03000000,
        32'h55020000,
        32'h03000000,
        32'h43020000,
        32'h03000000,
        32'h31020000,
        32'h03000000,
        32'h21020000,
        32'h03000000,
        32'h00000000,
        32'h00000000,
        32'h10000000,
        32'h11020000,
        32'h03000000,
        32'h612e3030,
        32'h6970672d,
        32'h786e6c78,
        32'h15000000,
        32'h02000000,
        32'h04000000,
        32'h00000030,
        32'h30303440,
        32'h01000000,
        32'h00800000,
        32'h00000030,
        32'h67000000,
        32'h03000000,
        32'h023e1800,
        32'h06000000,
        32'h00000000,
        32'h52010000,
        32'h03000000,
        32'h41010000,
        32'h03000000,
        32'h7774656e,
        32'h08000000,
        32'h00687465,
        32'h72776f6c,
        32'h0c000000,
        32'h00000000,
        32'h30303033,
        32'h2d637369,
        32'h01000000,
        32'h02000000,
        32'h00000000,
        32'he40c0000,
        32'hd9010000,
        32'h03000000,
        32'hc7010000,
        32'h03000000,
        32'h67000000,
        32'h03000000,
        32'h746f6c73,
        32'h2d636d6d,
        32'h0d000000,
        32'h00000030,
        32'h01000000,
        32'hb8010000,
        32'h03000000,
        32'ha1010000,
        32'h03000000,
        32'h90010000,
        32'h03000000,
        32'h80010000,
        32'h03000000,
        32'h746e696b,
        32'h08000000,
        32'h00100000,
        32'h00000020,
        32'h67000000,
        32'h03000000,
        32'h02000000,
        32'h08000000,
        32'h03000000,
        32'h04000000,
        32'h00000000,
        32'h04000000,
        32'h01000000,
        32'h04000000,
        32'h00612e30,
        32'h6970732d,
        32'h786e6c78,
        32'h302e322d,
        32'h7370782c,
        32'h1b000000,
        32'h03000000,
        32'h30303030,
        32'h40697073,
        32'h01000000,
        32'h04000000,
        32'h04000000,
        32'h02000000,
        32'h04000000,
        32'h01000000,
        32'h04000000,
        32'h03000000,
        32'h04000000,
        32'h00c20100,
        32'h04000000,
        32'h80f0fa02,
        32'h04000000,
        32'h00100000,
        32'h00000010,
        32'h67000000,
        32'h03000000,
        32'h3631736e,
        32'h08000000,
        32'h00000030,
        32'h30303140,
        32'h01000000,
        32'h006c6f72,
        32'h0b010000,
        32'h03000000,
        32'h00000000,
        32'h00000000,
        32'h10000000,
        32'hffff0000,
        32'hf7000000,
        32'h03000000,
        32'h2d677562,
        32'h63736972,
        32'h10000000,
        32'h00003040,
        32'h6f72746e,
        32'h75626564,
        32'h02000000,
        32'hb5000000,
        32'h03000000,
        32'h28010000,
        32'h03000000,
        32'h15010000,
        32'h03000000,
        32'h00000000,
        32'h00000000,
        32'h10000000,
        32'h09000000,
        32'h0b000000,
        32'hf7000000,
        32'h03000000,
        32'h00000000,
        32'h00306369,
        32'h63736972,
        32'h0c000000,
        32'h01000000,
        32'h04000000,
        32'h00000000,
        32'h04000000,
        32'h00000000,
        32'h30306340,
        32'h6f72746e,
        32'h70757272,
        32'h01000000,
        32'h006c6f72,
        32'h0b010000,
        32'h03000000,
        32'h00000000,
        32'h00000000,
        32'h10000000,
        32'h07000000,
        32'h03000000,
        32'hf7000000,
        32'h03000000,
        32'h30746e69,
        32'h63736972,
        32'h0d000000,
        32'h00000030,
        32'h30324074,
        32'h01000000,
        32'h00000000,
        32'h00007375,
        32'h706d6973,
        32'h2d657261,
        32'h61697261,
        32'h1b000000,
        32'h03000000,
        32'h0f000000,
        32'h03000000,
        32'h00000000,
        32'h03000000,
        32'h01000000,
        32'h02000000,
        32'h00000000,
        32'h00000074,
        32'h72616568,
        32'h0a000000,
        32'h00000000,
        32'h01000000,
        32'h0c000000,
        32'h00000064,
        32'h61656274,
        32'h01000000,
        32'h64656c2d,
        32'h1b000000,
        32'h03000000,
        32'h7364656c,
        32'h02000000,
        32'h00000000,
        32'h00000000,
        32'h10000000,
        32'h00007972,
        32'h5b000000,
        32'h03000000,
        32'h30303030,
        32'h6f6d656d,
        32'h02000000,
        32'h02000000,
        32'hb5000000,
        32'h03000000,
        32'h6e692d75,
        32'h63736972,
        32'h0f000000,
        32'ha0000000,
        32'h03000000,
        32'h8f000000,
        32'h03000000,
        32'h72656c6c,
        32'h6f632d74,
        32'h65746e69,
        32'h85000000,
        32'h03000000,
        32'h76732c76,
        32'h7c000000,
        32'h03000000,
        32'h66616d69,
        32'h72000000,
        32'h03000000,
        32'h63736972,
        32'h69726120,
        32'h1b000000,
        32'h03000000,
        32'h79616b6f,
        32'h05000000,
        32'h00000000,
        32'h04000000,
        32'h00757063,
        32'h04000000,
        32'h80f0fa02,
        32'h04000000,
        32'h00000030,
        32'h01000000,
        32'h38000000,
        32'h03000000,
        32'h0f000000,
        32'h03000000,
        32'h00000000,
        32'h03000000,
        32'h73757063,
        32'h02000000,
        32'h30323531,
        32'h30303030,
        32'h7261752f,
        32'h2c000000,
        32'h03000000,
        32'h736f6863,
        32'h00657261,
        32'h61697261,
        32'h26000000,
        32'h03000000,
        32'h2d657261,
        32'h61697261,
        32'h1b000000,
        32'h03000000,
        32'h0f000000,
        32'h03000000,
        32'h00000000,
        32'h03000000,
        32'h01000000,
        32'h00000000,
        32'h00000000,
        32'hd2020000,
        32'h10000000,
        32'h28000000,
        32'h38000000,
        32'hedfe0dd0,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h42413938,
        32'h33323130,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'ha0018402,
        32'h00000597,
        32'h0010041b,
        32'hf0ef057e,
        32'hebcff0ef,
        32'h00001517,
        32'he4060805,
        32'h85931141,
        32'h65f1b38d,
        32'h04450513,
        32'hbbd9d9e5,
        32'h1517f78f,
        32'hefcff0ef,
        32'h00001517,
        32'he9450513,
        32'hbbfddc65,
        32'h1517fa0f,
        32'hf24ff0ef,
        32'h00001517,
        32'hebc50513,
        32'hc92984aa,
        32'h8556865e,
        32'hf4cff0ef,
        32'h00001517,
        32'h08090913,
        32'hf64ff0ef,
        32'h05130000,
        32'h1be383bf,
        32'h000a4503,
        32'h0bc50513,
        32'h80fff0ef,
        32'hf94ff0ef,
        32'h00001517,
        32'h00893503,
        32'h0c450513,
        32'h837ff0ef,
        32'h00093503,
        32'h0cc50513,
        32'hff2a1be3,
        32'h0a05000a,
        32'h8a13fdef,
        32'h05130000,
        32'h19e38b3f,
        32'h0007c503,
        32'h4a01ffef,
        32'h8d130ce5,
        32'h15178d3f,
        32'hf513817f,
        32'h05130000,
        32'h4cc11005,
        32'h09130801,
        32'h8b0ad33f,
        32'h46057101,
        32'h845ff0ef,
        32'h00001517,
        32'h4556857f,
        32'h05130000,
        32'hf0ef4546,
        32'h0dc50513,
        32'h8f7ff0ef,
        32'hf0ef0ce5,
        32'h1517909f,
        32'h88dff0ef,
        32'h00001517,
        32'h656289ff,
        32'h05130000,
        32'hf0ef4552,
        32'h0cc50513,
        32'h8ffff0ef,
        32'hf0ef0ce5,
        32'h1517911f,
        32'h8d5ff0ef,
        32'h00001517,
        32'h45228e7f,
        32'h05130000,
        32'hf0ef6502,
        32'h0d450513,
        32'h905ff0ef,
        32'h00001517,
        32'h915ff0ef,
        32'h00001517,
        32'h8526927f,
        32'h05130000,
        32'hf0ef0be5,
        32'h1517c905,
        32'he41ff0ef,
        32'h46057101,
        32'h0c450513,
        32'h80826125,
        32'h6c426be2,
        32'h7a4279e2,
        32'h64468526,
        32'h011354fd,
        32'h0cc50513,
        32'hc90ddeff,
        32'h8aaa1080,
        32'he862f05a,
        32'he0cae4a6,
        32'hf456e8a2,
        32'h54798082,
        32'h6b4a6aea,
        32'h794a74ea,
        32'h8522547d,
        32'h0f450513,
        32'hc5dff0ef,
        32'hc65ff0ef,
        32'hc6dff0ef,
        32'hc75ff0ef,
        32'ha805c7ff,
        32'hf0ef4531,
        32'h4401f930,
        32'h849319fd,
        32'h15c50513,
        32'he7990369,
        32'h1c639041,
        32'h8c49cb7f,
        32'h03051413,
        32'hcc5ff0ef,
        32'h04040413,
        32'h892af15f,
        32'h854a0007,
        32'h07b30400,
        32'hc69ff0ef,
        32'h05938622,
        32'h1ee3cfff,
        32'h84133e80,
        32'h0a93e951,
        32'hd1dff0ef,
        32'h0ff67613,
        32'h0015161b,
        32'h0ff47593,
        32'h0ff5f593,
        32'hf61ff0ef,
        32'h0104559b,
        32'h45010184,
        32'h9be30785,
        32'h00f106b3,
        32'h567d4781,
        32'h842e84aa,
        32'hed56f152,
        32'hfd26e1a2,
        32'hf54e7155,
        32'h15428d3d,
        32'h979b1701,
        32'hd79b0105,
        32'h551b0105,
        32'h00c59513,
        32'h0045d51b,
        32'h15428d5d,
        32'h579b8082,
        32'h8d2d0045,
        32'h8d3d0045,
        32'hd79b8de9,
        32'h853e6402,
        32'he1114781,
        32'hc51157f9,
        32'hc91157fd,
        32'hfc6de07f,
        32'h4429b8ff,
        32'h05130000,
        32'hf0efe022,
        32'h80826105,
        32'h64a26442,
        32'h051bfc94,
        32'hf0efeb3f,
        32'h05130000,
        32'h842ae57f,
        32'h05134000,
        32'h0613fbdf,
        32'he822ec06,
        32'h80820141,
        32'h157d6402,
        32'h051bef3f,
        32'h051385a2,
        32'he8dff0ef,
        32'hf0efe022,
        32'h05134581,
        32'h11418082,
        32'h64a26442,
        32'h3513f565,
        32'h051b0124,
        32'h00f91b63,
        32'hecdff0ef,
        32'h842aed7f,
        32'heddff0ef,
        32'hee5ff0ef,
        32'hf0efe04a,
        32'hec064521,
        32'h08700613,
        32'h45018082,
        32'h64a26442,
        32'hf89ff0ef,
        32'h05130000,
        32'h15e3c00d,
        32'h892a347d,
        32'h45014581,
        32'h44857104,
        32'hec06e426,
        32'h1101ccff,
        32'h38450513,
        32'h60e26442,
        32'h852e65a2,
        32'h3cc50513,
        32'hcf5ff0ef,
        32'hf0efe42e,
        32'h05130000,
        32'he8221101,
        32'h64e27402,
        32'h147d0007,
        32'hd79b0185,
        32'hf0efeb5f,
        32'h06400413,
        32'hf0ef0ff4,
        32'hf0ef0ff5,
        32'h551bed5f,
        32'h75130104,
        32'hf0ef0184,
        32'hf0ef0404,
        32'hf0ef84aa,
        32'hf022e432,
        32'hf03ff06f,
        32'h8082557d,
        32'h00230785,
        32'h06c82683,
        32'h5178b77d,
        32'h00074703,
        32'h80824501,
        32'hdbb8577d,
        32'h02b6e163,
        32'h20000837,
        32'hfff58b85,
        32'h0737d3b8,
        32'h10600713,
        32'h00010320,
        32'h61630007,
        32'h200006b7,
        32'h200007b7,
        32'h10000793,
        32'h64a2d3b8,
        32'h644260e2,
        32'h577d2000,
        32'hf0ef4d65,
        32'h1517eb1f,
        32'h15024088,
        32'h4f450513,
        32'he3958b85,
        32'h57e0ff65,
        32'h849353f8,
        32'h07132000,
        32'h37fd0001,
        32'hd7a8dbb8,
        32'he822ec06,
        32'h1101e7ff,
        32'h52450513,
        32'h64a260e2,
        32'h4799e97f,
        32'h05130000,
        32'hf0ef9101,
        32'h2481eaff,
        32'h05130000,
        32'hd03c1660,
        32'hf0ef5765,
        32'h1517f51f,
        32'h02049513,
        32'hf0ef56e5,
        32'h15175064,
        32'h07932000,
        32'h37fd0001,
        32'h47292000,
        32'hf0efe426,
        32'h58e50513,
        32'h15178082,
        32'h8082c10c,
        32'h60e2ecff,
        32'h4503ed7f,
        32'h4503f55f,
        32'h002c1101,
        32'h694264e2,
        32'hfe9410e3,
        32'h00914503,
        32'h34610081,
        32'hf0ef0ff5,
        32'h00895533,
        32'h0413892a,
        32'hec26f022,
        32'h61456942,
        32'h70a2fe94,
        32'hf0ef0091,
        32'hf0ef3461,
        32'hfc3ff0ef,
        32'h002c0089,
        32'h4461892a,
        32'hec26f022,
        32'h00f58023,
        32'h00e580a3,
        32'h00074703,
        32'h771396e7,
        32'h1797b7f5,
        32'hf0ef8082,
        32'h60a2e509,
        32'h842ae406,
        32'h808200e7,
        32'h071300e7,
        32'h071300e7,
        32'h00a78223,
        32'h00e78023,
        32'h0ff57713,
        32'hf8000713,
        32'h100007b7,
        32'h0045959b,
        32'h0023dfe5,
        32'h01474783,
        32'h80820205,
        32'hc5031000,
        32'h00054503,
        32'h00238082,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h01f49493,
        32'hb8458593,
        32'hf1402573,
        32'h4009091b,
        32'h00448493,
        32'h0004a903,
        32'h00990933,
        32'hf1402973,
        32'hfe090ae3,
        32'h34402973,
        32'hff24c6e3,
        32'h02000937,
        32'h0124a023,
        32'h020004b7,
        32'h01a11113,
        32'h03249663,
        32'h00000493,
        32'h00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? {mem_H[addr_q],mem_L[addr_q]} : '0;
endmodule
