// COPYRIGHT HEADER


`ifndef __UVMT_CV32E40S_BASE_TEST_WORKAROUNDS_SV__
`define __UVMT_CV32E40S_BASE_TEST_WORKAROUNDS_SV__


// This file should be empty by the end of the project


`endif // __UVMT_CV32E40S_BASE_TEST_WORKAROUNDS_SV__
