`include "cv32e40p_asm_program_gen.sv"
