// COPYRIGHT HEADER


`ifndef __UVME_CV32_CONSTANTS_SV__
`define __UVME_CV32_CONSTANTS_SV__


parameter uvme_cv32_reset_default_clk_period = 10_000; // 10ns
parameter uvme_cv32_debug_default_clk_period = 10_000; // 10ns


`endif // __UVME_CV32_CONSTANTS_SV__
