// COPYRIGHT HEADER


`ifndef __UVML_HRTBT_TDEFS_SV__
`define __UVML_HRTBT_TDEFS_SV__





`endif // __UVML_HRTBT_TDEFS_SV__
