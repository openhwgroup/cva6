// Copyright 2024 Thales DIS France SAS
//
// Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.0
// You may obtain a copy of the License at https://solderpad.org/licenses/
//
// WT_NEW Cache Subsystem Adapter
// Bridges the WT_NEW cache (with privilege-level dual controllers) to the 
// standard CVA6 cache subsystem interface

module wt_new_cache_subsystem_adapter
  import ariane_pkg::*;
  import wt_cache_pkg::*;
  import wt_new_cache_pkg::*;
  import riscv::*;
  #(parameter config_pkg::cva6_cfg_t CVA6Cfg = config_pkg::cva6_cfg_empty,
    parameter type icache_areq_t = logic,
    parameter type icache_arsp_t = logic,
    parameter type icache_dreq_t = logic,
    parameter type icache_drsp_t = logic,
    parameter type dcache_req_i_t = logic,
    parameter type dcache_req_o_t = logic,
    parameter type icache_req_t = logic,
    parameter type icache_rtrn_t = logic,
    parameter int unsigned NumPorts = 4,
    parameter type noc_req_t = logic,
    parameter type noc_resp_t = logic)
   (
    input logic clk_i,
    input logic rst_ni,
    input riscv::priv_lvl_t priv_lvl_i,  // KEY: Privilege level for WT_NEW dual controllers
    
    // I$ interface (passthrough - WT_NEW only affects dcache)
    input logic icache_en_i,
    input logic icache_flush_i,
    output logic icache_miss_o,
    input icache_areq_t icache_areq_i,
    output icache_arsp_t icache_areq_o,
    input icache_dreq_t icache_dreq_i,
    output icache_drsp_t icache_dreq_o,
    
    // D$ interface (adapted to WT_NEW)
    input logic dcache_enable_i,
    input logic dcache_flush_i,
    output logic dcache_flush_ack_o,
    output logic dcache_miss_o,
    output logic [NumPorts-1:0][CVA6Cfg.DCACHE_SET_ASSOC-1:0] miss_vld_bits_o,
    input amo_req_t dcache_amo_req_i,
    output amo_resp_t dcache_amo_resp_o,
    input dcache_req_i_t [NumPorts-1:0] dcache_req_ports_i,
    output dcache_req_o_t [NumPorts-1:0] dcache_req_ports_o,
    output logic wbuffer_empty_o,
    output logic wbuffer_not_ni_o,
    
    // Memory interface
    output noc_req_t noc_req_o,
    input noc_resp_t noc_resp_i,
    input logic [63:0] inval_addr_i,
    input logic inval_valid_i,
    output logic inval_ready_o
   );

   // =========================================================================
   // ICACHE PASSTHROUGH - WT_NEW only affects DCACHE
   // =========================================================================
   
   // For now, use standard icache (WT_NEW is dcache innovation)
   cva6_icache #(
     .CVA6Cfg(CVA6Cfg),
     .icache_areq_t(icache_areq_t),
     .icache_arsp_t(icache_arsp_t),
     .icache_dreq_t(icache_dreq_t),
     .icache_drsp_t(icache_drsp_t),
     .icache_req_t(icache_req_t),
     .icache_rtrn_t(icache_rtrn_t)
   ) i_cva6_icache (
     .clk_i(clk_i),
     .rst_ni(rst_ni),
     .en_i(icache_en_i),
     .flush_i(icache_flush_i),
     .miss_o(icache_miss_o),
     .areq_i(icache_areq_i),
     .areq_o(icache_areq_o),
     .dreq_i(icache_dreq_i),
     .dreq_o(icache_dreq_o),
     .mem_rtrn_vld_i(1'b0),
     .mem_rtrn_i('0),
     .mem_data_req_o(),
     .mem_data_ack_i(1'b0),
     .mem_data_o()
   );

   // =========================================================================
   // WT_NEW DCACHE INTEGRATION
   // =========================================================================
   
`ifndef SYNTHESIS
   // Signal to indicate WT_NEW is active (visible in VCD)
   logic wt_new_cache_active;
   assign wt_new_cache_active = 1'b1;

   // Cache type override for VCD visibility
   logic [3:0] effective_dcache_type;
   assign effective_dcache_type = 4'd8; // WT_NEW value
`endif
   
   // =========================================================================
   // PRIVILEGE LEVEL MODIFIER FOR TESTING
   // =========================================================================
   
   // Modified privilege level for WT_NEW cache testing with performance optimization
   riscv::priv_lvl_t modified_priv_lvl;
   riscv::priv_lvl_t prev_priv_lvl;
   logic [31:0] priv_modifier_cycle_counter;
   logic priv_modifier_switch_event;
   logic priv_modifier_in_machine_mode;
   logic priv_modifier_in_user_mode;
   logic privilege_switch_detected;
   logic [3:0] switch_debounce_counter;
   
   // Instantiate privilege level modifier
   priv_lvl_modifier #(
     .SWITCH_PERIOD(100)  // Switch every 100 clock cycles
   ) i_priv_lvl_modifier (
     .clk_i(clk_i),
     .rst_ni(rst_ni),
     .actual_priv_lvl_i(priv_lvl_i),           // Actual privilege level (ignored)
     .modified_priv_lvl_o(modified_priv_lvl),  // Modified privilege level for testing
     .cycle_counter_o(priv_modifier_cycle_counter),
     .privilege_switch_event_o(priv_modifier_switch_event),
     .in_machine_mode_o(priv_modifier_in_machine_mode),
     .in_user_mode_o(priv_modifier_in_user_mode)
   );
   
   // =========================================================================
   // PRIVILEGE LEVEL SWITCHING PERFORMANCE OPTIMIZATION
   // =========================================================================
   
   // Track privilege level changes with debouncing for performance optimization
   always_ff @(posedge clk_i or negedge rst_ni) begin
     if (!rst_ni) begin
       prev_priv_lvl <= riscv::PRIV_LVL_M;
       privilege_switch_detected <= 1'b0;
       switch_debounce_counter <= '0;
     end else begin
       prev_priv_lvl <= modified_priv_lvl;
       
       // Detect privilege level switches with debouncing
       if (prev_priv_lvl != modified_priv_lvl) begin
         privilege_switch_detected <= 1'b1;
         switch_debounce_counter <= 4'd8; // 8-cycle debounce period
       end else if (switch_debounce_counter > 0) begin
         switch_debounce_counter <= switch_debounce_counter - 1;
       end else begin
         privilege_switch_detected <= 1'b0;
       end
     end
   end
   
   // Privilege level tracking for debugging with optimization hints
   riscv::priv_lvl_t current_priv_lvl;
   logic privilege_stable;
   
   assign current_priv_lvl = modified_priv_lvl; // Use modified privilege level
   assign privilege_stable = (switch_debounce_counter == 0) && !privilege_switch_detected;
   
   // Port arbitration - PROPER MULTI-PORT SUPPORT
   logic dcache_req_valid;
   logic [CVA6Cfg.PLEN-1:0] dcache_req_addr;
   logic dcache_req_we;
   logic [CVA6Cfg.DCACHE_LINE_WIDTH-1:0] dcache_req_wdata;
   logic [CVA6Cfg.DCACHE_LINE_WIDTH-1:0] dcache_resp_rdata;
   logic dcache_resp_hit;
   
   // AMO state machine type definition
   typedef enum logic [1:0] {
     AMO_IDLE,
     AMO_READ,
     AMO_MODIFY,
     AMO_WRITE
   } amo_state_t;
   
   // Forward declarations for AMO signals
   logic amo_req_valid;
   logic [63:0] amo_operand_a_q, amo_operand_b_q;
   logic [63:0] amo_result;
   amo_state_t amo_state_q;
   
   // Priority arbitration across all ports and AMO requests
   always_comb begin
     dcache_req_valid = 1'b0;
     dcache_req_addr  = '0;
     dcache_req_we    = 1'b0;
     dcache_req_wdata = '0;
     
     // AMO requests have highest priority
     if (amo_req_valid) begin
       dcache_req_valid = 1'b1;
       dcache_req_addr  = amo_operand_a_q[CVA6Cfg.PLEN-1:0];
       if (amo_state_q == AMO_WRITE) begin
         dcache_req_we = 1'b1;
         dcache_req_wdata = {{CVA6Cfg.DCACHE_LINE_WIDTH-64{1'b0}}, amo_result};
       end else begin
         dcache_req_we = 1'b0;
         dcache_req_wdata = '0;
       end
     end else begin
       // Regular port arbitration - port 0 has highest priority
       for (int i = NumPorts-1; i >= 0; i--) begin
         if (dcache_req_ports_i[i].data_req) begin
           dcache_req_valid = 1'b1;
           dcache_req_addr  = {{CVA6Cfg.PLEN-CVA6Cfg.XLEN{1'b0}}, dcache_req_ports_i[i].address_tag, dcache_req_ports_i[i].address_index};
           dcache_req_we    = dcache_req_ports_i[i].data_we;
           dcache_req_wdata = {{CVA6Cfg.DCACHE_LINE_WIDTH-CVA6Cfg.XLEN{1'b0}}, dcache_req_ports_i[i].data_wdata};
         end
       end
     end
   end
   
   // Performance counters for WT_NEW cache
   logic [63:0] wt_new_hit_count, wt_new_miss_count, wt_new_switch_count;
   
   // Dummy signals for debug outputs
   priv_lvl_t dummy_effective_priv;
   logic dummy_priv_override;
   logic [31:0] dummy_cycle_counter;
   
   // Instantiate the actual WT_NEW cache with modified privilege level
   wt_new_cache_subsystem #(
     .CVA6Cfg(CVA6Cfg),
     .NUM_DUAL_SETS(wt_new_cache_pkg::NUM_DUAL_SETS),
     .axi_req_t(noc_req_t),
     .axi_rsp_t(noc_resp_t)
   ) i_wt_new_cache (
     .clk_i(clk_i),
     .rst_ni(rst_ni),
     .priv_lvl_i(modified_priv_lvl),  // Use modified privilege level for predictable switching
     
     // NEW: Test mode control
     .test_mode_enable_i(1'b0),  // Default to real mode
     
     // Cache interface
     .req_i(dcache_req_valid & dcache_enable_i),
     .addr_i(dcache_req_addr),
     .we_i(dcache_req_we),
     .wdata_i(dcache_req_wdata),
     .rdata_o(dcache_resp_rdata),
     .hit_o(dcache_resp_hit),
     
     // Memory interface for miss handling
     .axi_data_req_o(noc_req_o),
     .axi_data_rsp_i(noc_resp_i),
     
     // Performance monitoring
     .hit_count_o(wt_new_hit_count),
     .miss_count_o(wt_new_miss_count),
     .switch_count_o(wt_new_switch_count),
     
     // NEW: Debug outputs for privilege mode control
     .effective_priv_lvl_o(dummy_effective_priv),
     .priv_mode_override_o(dummy_priv_override),
     .test_cycle_counter_o(dummy_cycle_counter)
   );
   
   // Map responses back to ports - PROPER CACHE BEHAVIOR with blocking on misses!
   always_comb begin
     // Initialize all ports
     for (int i = 0; i < NumPorts; i++) begin
       dcache_req_ports_o[i] = '0;
     end
     
     // Handle all port requests with proper cache blocking behavior
     for (int i = 0; i < NumPorts; i++) begin
       if (dcache_req_ports_i[i].data_req) begin
         // Grant immediately for all requests
         dcache_req_ports_o[i].data_gnt = 1'b1;
         
         // Handle kill requests immediately - this is critical for load unit
         if (dcache_req_ports_i[i].kill_req) begin
           dcache_req_ports_o[i].data_rvalid = 1'b1; // Acknowledge kill immediately
           dcache_req_ports_o[i].data_rdata  = '0;   // No data for killed requests
           dcache_req_ports_o[i].data_ruser  = '0;   // No user data for killed requests
           dcache_req_ports_o[i].data_rid    = dcache_req_ports_i[i].data_id; // Echo back ID
         end else begin
           // PROPER CACHE BEHAVIOR: Only respond when cache has valid data
           if (dcache_resp_hit) begin
             // Cache hit - respond immediately with valid data
             dcache_req_ports_o[i].data_rvalid = 1'b1;
             dcache_req_ports_o[i].data_rdata  = dcache_resp_rdata[CVA6Cfg.XLEN-1:0];
             dcache_req_ports_o[i].data_ruser  = '0;
             dcache_req_ports_o[i].data_rid    = dcache_req_ports_i[i].data_id;
           end else begin
             // Cache miss - DO NOT respond until cache completes memory fetch
             // This allows the cache miss handling FSM to work properly
             dcache_req_ports_o[i].data_rvalid = 1'b0; // Block until cache ready
             dcache_req_ports_o[i].data_rdata  = '0;
             dcache_req_ports_o[i].data_ruser  = '0;
             dcache_req_ports_o[i].data_rid    = dcache_req_ports_i[i].data_id;
           end
         end
       end
     end
   end
   
   // =========================================================================
   // CACHE MISS TRACKING (Cache handles its own memory interface)
   // =========================================================================
   
   // Simple cache miss detection for monitoring
   logic cache_miss;
   assign cache_miss = dcache_req_valid & ~dcache_resp_hit;
   
   // =========================================================================
   // CACHE FLUSH MECHANISM
   // =========================================================================
   
   // Flush state machine for proper cache invalidation
   typedef enum logic [1:0] {
     FLUSH_IDLE,
     FLUSH_ACTIVE,
     FLUSH_WAIT_COMPLETE
   } flush_state_t;
   
   flush_state_t flush_state_q, flush_state_d;
   logic [31:0] flush_counter;
   logic flush_complete;
   
   always_ff @(posedge clk_i or negedge rst_ni) begin
     if (!rst_ni) begin
       flush_state_q <= FLUSH_IDLE;
       flush_counter <= '0;
     end else begin
       flush_state_q <= flush_state_d;
       
       if (flush_state_q == FLUSH_ACTIVE) begin
         flush_counter <= flush_counter + 1;
       end else begin
         flush_counter <= '0;
       end
     end
   end
   
   always_comb begin
     flush_state_d = flush_state_q;
     flush_complete = 1'b0;
     
     case (flush_state_q)
       FLUSH_IDLE: begin
         if (dcache_flush_i) begin
           flush_state_d = FLUSH_ACTIVE;
         end
       end
       FLUSH_ACTIVE: begin
         // Allow time for cache flush operations
         if (flush_counter >= 16) begin // Give enough cycles for cache invalidation
           flush_state_d = FLUSH_WAIT_COMPLETE;
           flush_complete = 1'b1;
         end
       end
       FLUSH_WAIT_COMPLETE: begin
         flush_complete = 1'b1;
         if (!dcache_flush_i) begin
           flush_state_d = FLUSH_IDLE;
         end
       end
       default: begin
         flush_state_d = FLUSH_IDLE;
         flush_complete = 1'b0;
       end
     endcase
   end

   // Cache control signals
   assign dcache_flush_ack_o = flush_complete;
   assign dcache_miss_o = cache_miss;
   
   // =========================================================================
   // PERFORMANCE COUNTER SUPPORT - miss_vld_bits tracking
   // =========================================================================
   
   // Track cache misses for performance counters
   logic [NumPorts-1:0][CVA6Cfg.DCACHE_SET_ASSOC-1:0] miss_vld_bits;
   
   always_comb begin
     miss_vld_bits = '0;
     
     // Track misses per port
     for (int i = 0; i < NumPorts; i++) begin
       if (dcache_req_ports_i[i].data_req && ~dcache_resp_hit) begin
         // For WT_NEW cache, we can track misses in way 0 for simplicity
         // This gives visibility into cache miss patterns per port
         miss_vld_bits[i][0] = 1'b1;
       end
     end
   end
   
   assign miss_vld_bits_o = miss_vld_bits;
   
   // =========================================================================
   // AMO (Atomic Memory Operations) SUPPORT
   // =========================================================================
   
   // AMO state machine for atomic operations
   amo_state_t amo_state_d;
   logic [1:0] amo_size_q;
   amo_t amo_op_q;
   logic [63:0] amo_read_data;
   
   // Register AMO request
   always_ff @(posedge clk_i or negedge rst_ni) begin
     if (!rst_ni) begin
       amo_state_q <= AMO_IDLE;
       amo_operand_a_q <= '0;
       amo_operand_b_q <= '0;
       amo_size_q <= '0;
       amo_op_q <= AMO_NONE;
       amo_read_data <= '0;
     end else begin
       amo_state_q <= amo_state_d;
       
       // Capture AMO request
       if (dcache_amo_req_i.req && amo_state_q == AMO_IDLE) begin
         amo_operand_a_q <= dcache_amo_req_i.operand_a;
         amo_operand_b_q <= dcache_amo_req_i.operand_b;
         amo_size_q <= dcache_amo_req_i.size;
         amo_op_q <= dcache_amo_req_i.amo_op;
       end
       
       // Capture read data during AMO_READ state
       if (amo_state_q == AMO_READ && dcache_resp_hit) begin
         amo_read_data <= dcache_resp_rdata;
       end
     end
   end
   
   // AMO operation logic
   always_comb begin
     amo_result = amo_read_data; // Default to read data
     
     case (amo_op_q)
       AMO_SWAP: amo_result = amo_operand_b_q;
       AMO_ADD:  amo_result = amo_read_data + amo_operand_b_q;
       AMO_AND:  amo_result = amo_read_data & amo_operand_b_q;
       AMO_OR:   amo_result = amo_read_data | amo_operand_b_q;
       AMO_XOR:  amo_result = amo_read_data ^ amo_operand_b_q;
       AMO_MAX:  amo_result = ($signed(amo_read_data) > $signed(amo_operand_b_q)) ? amo_read_data : amo_operand_b_q;
       AMO_MIN:  amo_result = ($signed(amo_read_data) < $signed(amo_operand_b_q)) ? amo_read_data : amo_operand_b_q;
       AMO_MAXU: amo_result = (amo_read_data > amo_operand_b_q) ? amo_read_data : amo_operand_b_q;
       AMO_MINU: amo_result = (amo_read_data < amo_operand_b_q) ? amo_read_data : amo_operand_b_q;
       default:  amo_result = amo_read_data;
     endcase
   end
   
   // AMO state machine
   always_comb begin
     amo_state_d = amo_state_q;
     amo_req_valid = 1'b0;
     
     case (amo_state_q)
       AMO_IDLE: begin
         if (dcache_amo_req_i.req) begin
           amo_state_d = AMO_READ;
         end
       end
       AMO_READ: begin
         amo_req_valid = 1'b1; // Generate read request
         if (dcache_resp_hit) begin
           amo_state_d = AMO_MODIFY;
         end
       end
       AMO_MODIFY: begin
         // Computation happens combinatorially
         amo_state_d = AMO_WRITE;
       end
       AMO_WRITE: begin
         amo_req_valid = 1'b1; // Generate write request
         if (dcache_resp_hit) begin
           amo_state_d = AMO_IDLE;
         end
       end
     endcase
   end
   
   // AMO response generation
   always_comb begin
     dcache_amo_resp_o.ack = 1'b0;
     dcache_amo_resp_o.result = '0;
     
     if (amo_state_q == AMO_WRITE && dcache_resp_hit) begin
       dcache_amo_resp_o.ack = 1'b1;
       // Return original read data for most AMOs, result for SWAP
       dcache_amo_resp_o.result = (amo_op_q == AMO_SWAP) ? amo_result : amo_read_data;
     end
   end
   
   // Write buffer (WT_NEW is write-through, so always empty)
   assign wbuffer_empty_o = 1'b1;
   assign wbuffer_not_ni_o = 1'b0;
   
   // Invalidation interface
   assign inval_ready_o = 1'b1;

endmodule
