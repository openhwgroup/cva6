/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 835;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h0a0d2165_6e6f6420,
        64'h00000000_00206567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f63,
        64'h00000000_00000009,
        64'h3a656d61_6e090a0d,
        64'h00093a73_65747562,
        64'h69727474_61090a0d,
        64'h00000009_3a61626c,
        64'h20747361_6c090a0d,
        64'h0000093a_61626c20,
        64'h74737269_66090a0d,
        64'h00000000_00000000,
        64'h09202020_20203a64,
        64'h69756720_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_00000000,
        64'h093a6469_75672065,
        64'h70797420_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20747067,
        64'h00000009_20203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20657a69_73090a0d,
        64'h00000009_3a736569,
        64'h72746e65_206e6f69,
        64'h74697472_61702072,
        64'h65626d75_6e090a0d,
        64'h00000009_2020203a,
        64'h61626c20_73656972,
        64'h746e6520_6e6f6974,
        64'h69747261_70090a0d,
        64'h00093a61_646c2070,
        64'h756b6361_62090a0d,
        64'h00000000_00000000,
        64'h093a6162_6c20746e,
        64'h65727275_63090a0d,
        64'h00000009_3a646576,
        64'h72657365_72090a0d,
        64'h00093a72_65646165,
        64'h685f6372_63090a0d,
        64'h00000000_00000909,
        64'h3a657a69_73090a0d,
        64'h00000009_3a6e6f69,
        64'h73697665_72090a0d,
        64'h0000093a_65727574,
        64'h616e6769_73090a0d,
        64'h00000000_003a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20747067,
        64'h0000203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_63206473,
        64'h00000000_0000000a,
        64'h0d216465_7a696c61,
        64'h6974696e_69206473,
        64'h00000000_0a0d676e,
        64'h69746978_65202e2e,
        64'h2e647320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f63,
        64'h00000000_0000002e,
        64'h0000000a_0d202e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e69,
        64'h00000031_34646d63,
        64'h00000035_35646d63,
        64'h00000000_30646d63,
        64'h00000020_3a206573,
        64'h6e6f7073_65720920,
        64'h00000000_0020646e,
        64'h616d6d6f_63204453,
        64'h00000000_00000a0d,
        64'h65736e6f_70736572,
        64'h20647320_64696c61,
        64'h7620646e_69662074,
        64'h6f6e2064_6c756f63,
        64'h00000000_203f3f79,
        64'h74706d65_20746f6e,
        64'h206f6669_66207872,
        64'h00000000_00000a0d,
        64'h2164657a_696c6169,
        64'h74696e69_20495053,
        64'h00000000_00007830,
        64'h203a7375_74617473,
        64'h00000000_00000a0d,
        64'h49505320_74696e69,
        64'h00000a0d_21646c72,
        64'h6f57206f_6c6c6548,
        64'h00000000_00006564,
        64'h6f6d2d79_6870006f,
        64'h69646d2d_7361682c,
        64'h786e6c78_006c616e,
        64'h7265746e_692d6573,
        64'h752c786e_6c780067,
        64'h6e6f702d_676e6970,
        64'h2d78742c_786e6c78,
        64'h00687464_69772d64,
        64'h692d6978_612d732c,
        64'h786e6c78_00676e6f,
        64'h702d676e_69702d78,
        64'h722c786e_6c780065,
        64'h636e6174_736e692c,
        64'h786e6c78_006f6964,
        64'h6d2d6564_756c636e,
        64'h692c786e_6c78006b,
        64'h63616270_6f6f6c2d,
        64'h6c616e72_65746e69,
        64'h2d656475_6c636e69,
        64'h2c786e6c_78007372,
        64'h65666675_622d6c61,
        64'h626f6c67_2d656475,
        64'h6c636e69_2c786e6c,
        64'h78007865_6c707564,
        64'h2c786e6c_7800656c,
        64'h646e6168_2d796870,
        64'h00737365_72646461,
        64'h2d63616d_2d6c6163,
        64'h6f6c0070_772d656c,
        64'h62617369_64007365,
        64'h676e6172_2d656761,
        64'h746c6f76_0079636e,
        64'h65757165_72662d78,
        64'h616d2d69_7073006f,
        64'h69746172_2d6b6373,
        64'h2c786e6c_78007374,
        64'h69622d72_6566736e,
        64'h6172742d_6d756e2c,
        64'h786e6c78_00737469,
        64'h622d7373_2d6d756e,
        64'h2c786e6c_78007473,
        64'h6978652d_6f666966,
        64'h2c786e6c_7800796c,
        64'h696d6166_2c786e6c,
        64'h78006874_6469772d,
        64'h6f692d67_65720074,
        64'h66696873_2d676572,
        64'h00737470_75727265,
        64'h746e6900_746e6572,
        64'h61702d74_70757272,
        64'h65746e69_00646565,
        64'h70732d74_6e657272,
        64'h75630076_65646e2c,
        64'h76637369_72007974,
        64'h69726f69_72702d78,
        64'h616d2c76_63736972,
        64'h0073656d_616e2d67,
        64'h65720064_65646e65,
        64'h7478652d_73747075,
        64'h72726574_6e690073,
        64'h65676e61_7200656c,
        64'h646e6168_702c7875,
        64'h6e696c00_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h02000000_02000000,
        64'h03000000_bb000000,
        64'h04000000_03000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h01000000_67000000,
        64'h04000000_03000000,
        64'h00000000_7968702d,
        64'h74656e72_65687465,
        64'h5b000000_0d000000,
        64'h03000000_00000000,
        64'h35313963_2e633130,
        64'h3064692d_7968702d,
        64'h74656e72_65687465,
        64'h1b000000_19000000,
        64'h03000000_00003040,
        64'h7968702d_74656e72,
        64'h65687465_01000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_6f69646d,
        64'h01000000_00000000,
        64'h64692d69_696d6772,
        64'ha2020000_09000000,
        64'h03000000_01000000,
        64'h94020000_04000000,
        64'h03000000_00000000,
        64'h82020000_04000000,
        64'h03000000_01000000,
        64'h70020000_04000000,
        64'h03000000_04000000,
        64'h5c020000_04000000,
        64'h03000000_01000000,
        64'h4a020000_04000000,
        64'h03000000_00657469,
        64'h6c74656e_72656874,
        64'h655f6978_615f786e,
        64'h6c785f69_3c020000,
        64'h18000000_03000000,
        64'h01000000_2a020000,
        64'h04000000_03000000,
        64'h00000000_0b020000,
        64'h04000000_03000000,
        64'h01000000_ef010000,
        64'h04000000_03000000,
        64'h01000000_e3010000,
        64'h04000000_03000000,
        64'h00000100_00000000,
        64'h00000030_00000000,
        64'h67000000_10000000,
        64'h03000000_03000000,
        64'hd8010000_04000000,
        64'h03000000_00002201,
        64'h00350a00_c6010000,
        64'h06000000_03000000,
        64'h00000000_03000000,
        64'h25010000_08000000,
        64'h03000000_02000000,
        64'h14010000_04000000,
        64'h03000000_006b726f,
        64'h7774656e_5b000000,
        64'h08000000_03000000,
        64'h0000612e_30302e31,
        64'h2d657469_6c74656e,
        64'h72656874_652d7370,
        64'h782c786e_6c780030,
        64'h2e332d65_74696c74,
        64'h656e7265_6874652d,
        64'h6978612c_786e6c78,
        64'h1b000000_37000000,
        64'h03000000_00000030,
        64'h30303030_30303340,
        64'h74656e72_65687465,
        64'h01000000_02000000,
        64'h02000000_bb010000,
        64'h00000000_03000000,
        64'he40c0000_e40c0000,
        64'hac010000_08000000,
        64'h03000000_20bcbe00,
        64'h9a010000_04000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00000000,
        64'h746f6c73_2d697073,
        64'h2d636d6d_1b000000,
        64'h0d000000_03000000,
        64'h00000030_40636d6d,
        64'h01000000_04000000,
        64'h8b010000_04000000,
        64'h03000000_08000000,
        64'h74010000_04000000,
        64'h03000000_01000000,
        64'h63010000_04000000,
        64'h03000000_01000000,
        64'h53010000_04000000,
        64'h03000000_00377865,
        64'h746e696b_47010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000020_00000000,
        64'h67000000_10000000,
        64'h03000000_02000000,
        64'h02000000_25010000,
        64'h08000000_03000000,
        64'h02000000_14010000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00612e30_302e322d,
        64'h6970732d_7370782c,
        64'h786e6c78_00622e30,
        64'h302e322d_6970732d,
        64'h7370782c_786e6c78,
        64'h1b000000_28000000,
        64'h03000000_00000000,
        64'h30303030_30303032,
        64'h40697073_2d737078,
        64'h01000000_02000000,
        64'h04000000_3a010000,
        64'h04000000_03000000,
        64'h02000000_30010000,
        64'h04000000_03000000,
        64'h01000000_25010000,
        64'h04000000_03000000,
        64'h02000000_14010000,
        64'h04000000_03000000,
        64'h00c20100_06010000,
        64'h04000000_03000000,
        64'h80f0fa02_4b000000,
        64'h04000000_03000000,
        64'h00100000_00000000,
        64'h00000010_00000000,
        64'h67000000_10000000,
        64'h03000000_00303537,
        64'h3631736e_1b000000,
        64'h08000000_03000000,
        64'h00000030_30303030,
        64'h30303140_74726175,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'hde000000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000000,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'hffff0000_01000000,
        64'hca000000_08000000,
        64'h03000000_00333130,
        64'h2d677562_65642c76,
        64'h63736972_1b000000,
        64'h10000000_03000000,
        64'h00003040_72656c6c,
        64'h6f72746e_6f632d67,
        64'h75626564_01000000,
        64'h02000000_02000000,
        64'hbb000000_04000000,
        64'h03000000_02000000,
        64'hb5000000_04000000,
        64'h03000000_03000000,
        64'hfb000000_04000000,
        64'h03000000_07000000,
        64'he8000000_04000000,
        64'h03000000_00000004,
        64'h00000000_0000000c,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h09000000_01000000,
        64'h0b000000_01000000,
        64'hca000000_10000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h00306369_6c702c76,
        64'h63736972_1b000000,
        64'h0c000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_00000000,
        64'h04000000_03000000,
        64'h00000000_30303030,
        64'h30306340_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'hde000000_08000000,
        64'h03000000_00000c00,
        64'h00000000_00000002,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h07000000_01000000,
        64'h03000000_01000000,
        64'hca000000_10000000,
        64'h03000000_00000000,
        64'h30746e69_6c632c76,
        64'h63736972_1b000000,
        64'h0d000000_03000000,
        64'h00000030_30303030,
        64'h30324074_6e696c63,
        64'h01000000_c3000000,
        64'h00000000_03000000,
        64'h00007375_622d656c,
        64'h706d6973_00636f73,
        64'h2d657261_622d656e,
        64'h61697261_2c687465,
        64'h1b000000_1f000000,
        64'h03000000_02000000,
        64'h0f000000_04000000,
        64'h03000000_02000000,
        64'h00000000_04000000,
        64'h03000000_00636f73,
        64'h01000000_02000000,
        64'h00000008_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h01000000_bb000000,
        64'h04000000_03000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00007573_63616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h10090000_ab020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h48090000_38000000,
        64'hf30b0000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_0000a001,
        64'h840202a5_85930000,
        64'h059701f4_14130010,
        64'h041bd5df_f0ef057e,
        64'h65a14505_f42ff0ef,
        64'hc4050513_00001517,
        64'hf1cff0ef_e4061141,
        64'hb375815a_f5aff0ef,
        64'hf3850513_00001517,
        64'hc61ff0ef_855e8662,
        64'h020aa583_f72ff0ef,
        64'hf3850513_00001517,
        64'hf59910e3_08048493,
        64'h080a0993_f8aff0ef,
        64'h2905cca5_05130000,
        64'h1517ff3a_1be3861f,
        64'hf0ef0a05_000a4503,
        64'hfa6ff0ef_f5c50513,
        64'h00001517_835ff0ef,
        64'h6888fb8f_f0eff5e5,
        64'h05130000_1517847f,
        64'hf0ef6488_fcaff0ef,
        64'hf6050513_00001517,
        64'h859ff0ef_fb898a13,
        64'h6088fe0f_f0eff665,
        64'h05130000_1517fe9a,
        64'h1be38b5f_f0ef0a05,
        64'h000a4503_f9098a13,
        64'hffeff0ef_f6450513,
        64'h00001517_ffaa19e3,
        64'h8d3ff0ef_0a050007,
        64'hc503014d_87b34a01,
        64'h81fff0ef_f8098d93,
        64'hf6850513_00001517,
        64'h8f3ff0ef_0ff97513,
        64'h837ff0ef_f6450513,
        64'h00001517_4c914d41,
        64'h020a8493_080a8993,
        64'h84fff0ef_d8c50513,
        64'h00001517_8ddff0ef,
        64'h8526861f_f0efe7e5,
        64'h05130000_1517c105,
        64'h84aa8a8a_d6dff0ef,
        64'h850a4605_710144ac,
        64'h87fff0ef_dbc50513,
        64'h00001517_8cdff0ef,
        64'h48e8891f_f0eff9e5,
        64'h05130000_15178dff,
        64'hf0ef48a8_8a3ff0ef,
        64'hf9050513_00001517,
        64'h931ff0ef_64a88b5f,
        64'hf0eff825_05130000,
        64'h1517943f_f0ef7088,
        64'h8c7ff0ef_f8450513,
        64'h00001517_955ff0ef,
        64'h6c888d9f_f0eff7e5,
        64'h05130000_1517927f,
        64'hf0ef48c8_8ebff0ef,
        64'hf8050513_00001517,
        64'h939ff0ef_48888fdf,
        64'hf0eff825_05130000,
        64'h151794bf_f0ef44c8,
        64'h90fff0ef_f8450513,
        64'h00001517_95dff0ef,
        64'h4488921f_f0eff865,
        64'h05130000_15179aff,
        64'hf0ef6088_933ff0ef,
        64'hf8850513_00001517,
        64'h93fff0ef_f7450513,
        64'h00001517_94bff0ef,
        64'he8850513_00001517,
        64'h9d9ff0ef_854e95df,
        64'hf0eff7a5_05130000,
        64'h1517c105_89aa848a,
        64'he69ff0ef_850a4585,
        64'h46057101_8b0a97df,
        64'hf0eff825_05130000,
        64'h1517892a_80826165,
        64'h6da26d42_6ce27c02,
        64'h7ba27b42_7ae26a06,
        64'h69a66946_64e67406,
        64'h70a6f904_01139adf,
        64'hf0eff8a5_05130000,
        64'h1517c905_e19ff0ef,
        64'h8c2e8baa_1880e46e,
        64'he86aec66_f85afc56,
        64'he0d2e4ce_e8caeca6,
        64'hf486f062_f45ef0a2,
        64'h7159bfe1_54798082,
        64'h61696baa_6b4a6aea,
        64'h7a0a79aa_794a74ea,
        64'h640e60ae_8522c7df,
        64'hf0efc89f_f0ef4531,
        64'h45814605_4401f890,
        64'h46e32009_091314fd,
        64'ha17ff0ef_fec50513,
        64'h00001517_e7990364,
        64'he7b30489_94639041,
        64'h29811442_8c49cb5f,
        64'hf0ef9041_03051413,
        64'h0085151b_cc3ff0ef,
        64'hfd241ae3_04040413,
        64'hff7a17e3_89aaf11f,
        64'hf0ef0a05_854e0007,
        64'hc5830144_07b30400,
        64'h0b934a01_c67ff0ef,
        64'h850a0400_05938622,
        64'h4981ff55_1ee3cfdf,
        64'hf0efe009_04133e80,
        64'h0b130fe0_0a932009,
        64'h09139081_1482bff5,
        64'hd17ff0ef_c501d25f,
        64'hf0ef4549_85a20ff6,
        64'h76130016_66130015,
        64'h161bf53f_f0ef0ff4,
        64'h7593f5bf_f0ef0ff5,
        64'hf5930084_559bf67f,
        64'hf0ef0ff5_f5930104,
        64'h559bf73f_f0ef4501,
        64'h0184559b_fee79be3,
        64'h078500c6_802300f1,
        64'h06b30800_0713567d,
        64'h4781842e_892ae55e,
        64'he95aed56_f152f54e,
        64'he58684b2_f94afd26,
        64'he1a27155_80829141,
        64'h15428d3d_8ff90057,
        64'h979b1701_67090107,
        64'hd79b0105_179b4105,
        64'h551b0105_151b8d2d,
        64'h00c59513_8da9893d,
        64'h0045d51b_8da99141,
        64'h15428d5d_05220085,
        64'h579b8082_07f57513,
        64'h8d2d0045_15938d2d,
        64'h8d3d0045_d51b0075,
        64'hd79b8de9_80820141,
        64'h853e6402_60a257f5,
        64'he1114781_f89ff0ef,
        64'hc51157f9_efbff0ef,
        64'hc91157fd_ec9ff0ef,
        64'hfc6de09f_f0ef347d,
        64'h4429b91f_f0ef14e5,
        64'h05130000_1517c8bf,
        64'hf0efe022_e4061141,
        64'h80826105_00153513,
        64'h64a26442_60e20004,
        64'h051bfc94_0ce3e3df,
        64'hf0efec5f_f0ef1765,
        64'h05130000_151785aa,
        64'h842ae59f_f0ef0290,
        64'h05134000_05b70770,
        64'h0613fbdf_f0ef4485,
        64'he822ec06_e4261101,
        64'h80820141_00153513,
        64'h157d6402_60a20004,
        64'h051bf05f_f0ef1b05,
        64'h051385a2_00001517,
        64'he8fff0ef_842ae9df,
        64'hf0efe022_e4060370,
        64'h05134581_06500613,
        64'h11418082_61056902,
        64'h64a26442_60e20015,
        64'h3513f565_05130004,
        64'h051b0124_986388bd,
        64'h00f91b63_45014785,
        64'hecfff0ef_ed3ff0ef,
        64'h842aed9f_f0ef84aa,
        64'hedfff0ef_ee3ff0ef,
        64'hee7ff0ef_892aef5f,
        64'hf0efe04a_e426e822,
        64'hec064521_1aa00593,
        64'h08700613_11018082,
        64'h61054505_64a26442,
        64'h60e2fe94_10e3f99f,
        64'hf0ef23c5_051385a2,
        64'h00001517_f23ff0ef,
        64'h842af31f_f0ef4501,
        64'h09500613_45814485,
        64'he822ec06_e4261101,
        64'hcbfff06f_61051fe5,
        64'h05130000_151760e2,
        64'h6442d95f_f0ef852e,
        64'h65a2cd9f_f0ef26e5,
        64'h05130000_1517ce5f,
        64'hf0ef8522_cebff0ef,
        64'he42eec06_27450513,
        64'h00001517_842ae822,
        64'h11018082_614564e2,
        64'h85267402_70a2d0df,
        64'hf0ef26a5_05130000,
        64'h1517f475_147d0007,
        64'hda6384aa_4187d79b,
        64'h0185179b_fabff0ef,
        64'heb5ff0ef_85320640,
        64'h04136622_ec1ff0ef,
        64'h0ff47513_ec9ff0ef,
        64'h0ff57513_0084551b,
        64'hed5ff0ef_0ff57513,
        64'h0104551b_ee1ff0ef,
        64'h0184551b_ee9ff0ef,
        64'h0404e513_febff0ef,
        64'h84aa842e_ec26f022,
        64'he432f406_7179f03f,
        64'hf06f0ff0_05138082,
        64'h557db7d9_00d70023,
        64'h078500f6_073306c8,
        64'h2683ff69_8b055178,
        64'hb77dd6b8_07850007,
        64'h470300f5_07338082,
        64'h4501d3b8_4719dbb8,
        64'h577d2000_07b702b6,
        64'he1630007_869b2000,
        64'h08372000_0537fff5,
        64'h8b85537c_20000737,
        64'hd3b82000_07b71060,
        64'h0713fff5_37fd0001,
        64'h03200793_04b76163,
        64'h0007871b_47812000,
        64'h06b7dbb8_57792000,
        64'h07b706b7_ee631000,
        64'h07938082_610564a2,
        64'hd3b84719_dbb86442,
        64'h60e20ff4_7513577d,
        64'h200007b7_e23ff0ef,
        64'h36050513_00001517,
        64'heb1ff0ef_91011502,
        64'h4088e39f_f0ef37e5,
        64'h05130000_1517e395,
        64'h8b852401_53fc57e0,
        64'hff658b05_06478493,
        64'h53f8d3b8_10600713,
        64'h200007b7_fff537fd,
        64'h00010640_0793d7a8,
        64'hdbb85779_e426e822,
        64'hec062000_07b71101,
        64'he7fff06f_61053ae5,
        64'h05130000_151764a2,
        64'h60e26442_d03c4799,
        64'he97ff0ef_3d450513,
        64'h00001517_f25ff0ef,
        64'h91010204_95132481,
        64'heafff0ef_3cc50513,
        64'h00001517_5064d03c,
        64'h16600793_ec3ff0ef,
        64'h40050513_00001517,
        64'hf51ff0ef_91010204,
        64'h95132481_edbff0ef,
        64'h3f850513_00001517,
        64'h5064d03c_10400793,
        64'h20000437_fff537fd,
        64'h000147a9_c3b84729,
        64'h200007b7_f03ff0ef,
        64'he426e822_ec064185,
        64'h05131101_00001517,
        64'h80822501_41088082,
        64'hc10c8082_610560e2,
        64'hee1ff0ef_00914503,
        64'hee9ff0ef_00814503,
        64'hf55ff0ef_ec06002c,
        64'h11018082_61456942,
        64'h64e27402_70a2fe94,
        64'h10e3f0bf_f0ef0091,
        64'h4503f13f_f0ef3461,
        64'h00814503_f81ff0ef,
        64'h0ff57513_002c0089,
        64'h553354e1_03800413,
        64'h892af406_e84aec26,
        64'hf0227179_80826145,
        64'h694264e2_740270a2,
        64'hfe9410e3_f4dff0ef,
        64'h00914503_f55ff0ef,
        64'h34610081_4503fc3f,
        64'hf0ef0ff5_7513002c,
        64'h0089553b_54e14461,
        64'h892af406_e84aec26,
        64'hf0227179_808200f5,
        64'h80230007_c78300e5,
        64'h80a397aa_81110007,
        64'h4703973e_00f57713,
        64'h88078793_00002797,
        64'hb7f50405_fa5ff0ef,
        64'h80820141_640260a2,
        64'he5090004_4503842a,
        64'he406e022_11418082,
        64'h00e78823_02000713,
        64'h00e78423_fc700713,
        64'h00e78623_470d0007,
        64'h822300e7_8023476d,
        64'h00e78623_f8000713,
        64'h00078223_100007b7,
        64'h808200a7_0023dfe5,
        64'h0207f793_01474783,
        64'h10000737_80820205,
        64'h75130147_c5031000,
        64'h07b78082_00054503,
        64'h808200b5_00238082,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_01f49493,
        64'h0010049b_9e458593,
        64'h00001597_f1402573,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'hfe091ee3_0004a903,
        64'h00092023_00990933,
        64'h00291913_f1402973,
        64'h020004b7_fe090ae3,
        64'h00897913_34402973,
        64'h10500073_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_0124a023,
        64'h00100913_020004b7,
        64'h1f5000ef_fec10113,
        64'h01000117_03249663,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
