// COPYRIGHT HEADER


`ifndef __UVME_CV32_REG_IGNORE_ALL_LIST_SV__
`define __UVME_CV32_REG_IGNORE_ALL_LIST_SV__


string  ignore_list = '{
   // TODO Add register blocks to CV32 ignore list for all RAL automated tests
   //      Ex: "block_name.reg_name", // One register at a time
   //      Ex: "block_name.*", // One block at a time
};


`endif // __UVME_${tb_name_uppercase}_REG_IGNORE_ALL_LIST_SV__
