// Copyright 2018 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.
//
// Author: Florian Zaruba, ETH Zurich
// Date: 15/04/2017
// Description: Top level testbench module. Instantiates the top level DUT, configures
//              the virtual interfaces and starts the test passed by +UVM_TEST+

`timescale 1ps/1ps

import ariane_pkg::*;
import uvm_pkg::*;

`include "uvm_macros.svh"

import "DPI-C" function read_elf(input string filename);
import "DPI-C" function byte get_section(output longint address, output longint len);
import "DPI-C" context function byte read_section(input longint address, inout byte buffer[]);

module ariane_tb;

    static uvm_cmdline_processor uvcl = uvm_cmdline_processor::get_inst();

    localparam int unsigned CLOCK_PERIOD = 20ns;
    // toggle with RTC period
    localparam int unsigned RTC_CLOCK_PERIOD = 30.517us;

    localparam NUM_WORDS = 2**25;
    logic clk_i;
    logic rst_ni;
    logic rtc_i;

    parameter  USE_HYPER_MODELS    = 1;

    wire [7:0]            w_hyper_dq0    ;
    wire [7:0]            w_hyper_dq1    ;
    wire                  w_hyper_ck     ;
    wire                  w_hyper_ckn    ;
    wire                  w_hyper_csn0   ;
    wire                  w_hyper_csn1   ;
    wire                  w_hyper_rwds0  ;
    wire                  w_hyper_rwds1  ;
    wire                  w_hyper_reset  ;

    wire [63:0]           w_gpios        ; 

    wire                  w_cva6_uart_rx ;
    wire                  w_cva6_uart_tx ;
   
    wire  [1:0] axi_hyper_cs_n_wire;
    wire        axi_hyper_ck_wire;
    wire        axi_hyper_ck_n_wire;
    wire        axi_hyper_rwds_o;
    wire        axi_hyper_rwds_i;
    wire        axi_hyper_rwds_oe;
    wire        axi_hyper_rwds_wire;
 
    wire  [7:0] axi_hyper_dq_i;
    wire  [7:0] axi_hyper_dq_o;
    wire        axi_hyper_dq_oe;
    wire  [7:0] axi_hyper_dq_wire;
 
    wire        axi_hyper_reset_n_wire;
    
    tristate_shim i_tristate_shim_rwds (
        .out_ena_i  (  axi_hyper_rwds_oe   ),
        .out_i      (  axi_hyper_rwds_o    ),
        .in_o       (  axi_hyper_rwds_i    ),
        .line_io    (  axi_hyper_rwds_wire )
    );
 
    for (genvar i = 0; i < 8; i++) begin
        tristate_shim i_tristate_shim_dq (
            .out_ena_i  ( axi_hyper_dq_oe       ),
            .out_i      ( axi_hyper_dq_o    [i] ),
            .in_o       ( axi_hyper_dq_i    [i] ),
            .line_io    ( axi_hyper_dq_wire [i] )
        );
    end
  
    longint unsigned cycles;
    longint unsigned max_cycles;

    logic [31:0] exit_o;

    string binary = "";

    genvar j;
    generate
       for (j=0; j<32; j++) begin
          assign w_gpios[63-j] = w_gpios[j] ? 1 : 0 ;          
        end
    endgenerate

    al_saqr #(
        .NUM_WORDS         ( NUM_WORDS ),
        .InclSimDTM        ( 1'b1      ),
        .StallRandomOutput ( 1'b1      ),
        .StallRandomInput  ( 1'b1      )
    ) dut (
        .clk_i,
        .rst_ni,
        .rtc_i,
        .exit_o,
        .pad_hyper_dq0       ( w_hyper_dq0            ),
        .pad_hyper_dq1       ( w_hyper_dq1            ),
        .pad_hyper_ck        ( w_hyper_ck             ),
        .pad_hyper_ckn       ( w_hyper_ckn            ),
        .pad_hyper_csn0      ( w_hyper_csn0           ),
        .pad_hyper_csn1      ( w_hyper_csn1           ),
        .pad_hyper_rwds0     ( w_hyper_rwds0          ),
        .pad_hyper_rwds1     ( w_hyper_rwds1          ),
        .pad_hyper_reset     ( w_hyper_reset          ),
        .pad_gpio            ( w_gpios                ),
        .cva6_uart_rx_i      ( w_cva6_uart_rx         ),
        .cva6_uart_tx_o      ( w_cva6_uart_tx         ),
        .axi_hyper_cs_no     ( axi_hyper_cs_n_wire    ),
        .axi_hyper_ck_o      ( axi_hyper_ck_wire      ),
        .axi_hyper_ck_no     ( axi_hyper_ck_n_wire    ),
        .axi_hyper_rwds_o    ( axi_hyper_rwds_o       ),
        .axi_hyper_rwds_i    ( axi_hyper_rwds_i       ),
        .axi_hyper_rwds_oe_o ( axi_hyper_rwds_oe      ),
        .axi_hyper_dq_i      ( axi_hyper_dq_i         ),
        .axi_hyper_dq_o      ( axi_hyper_dq_o         ),
        .axi_hyper_dq_oe_o   ( axi_hyper_dq_oe        ),
        .axi_hyper_reset_no  ( axi_hyper_reset_n_wire )
   );

   s27ks0641 #(
         /*.mem_file_name ( "s27ks0641.mem"    ),*/
         .TimingModel   ( "S27KS0641DPBHI020"    )
     ) i_s27ks0641 (
       .DQ7           ( axi_hyper_dq_wire[7]      ),
       .DQ6           ( axi_hyper_dq_wire[6]      ),
       .DQ5           ( axi_hyper_dq_wire[5]      ),
       .DQ4           ( axi_hyper_dq_wire[4]      ),
       .DQ3           ( axi_hyper_dq_wire[3]      ),
       .DQ2           ( axi_hyper_dq_wire[2]      ),
       .DQ1           ( axi_hyper_dq_wire[1]      ),
       .DQ0           ( axi_hyper_dq_wire[0]      ),
       .RWDS          ( axi_hyper_rwds_wire       ),
       .CSNeg         ( axi_hyper_cs_n_wire[0]    ),
       .CK            ( axi_hyper_ck_wire         ),
       .CKNeg         ( axi_hyper_ck_n_wire       ),
       .RESETNeg      ( axi_hyper_reset_n_wire    )
     );

// Hyperram and hyperflash modules
   generate
      if(USE_HYPER_MODELS == 1) begin
         s27ks0641 #(
            .TimingModel  ("S27KS0641DPBHI020")
         ) hyperram_model (
            .DQ7      ( w_hyper_dq0[7] ),
            .DQ6      ( w_hyper_dq0[6] ),
            .DQ5      ( w_hyper_dq0[5] ),
            .DQ4      ( w_hyper_dq0[4] ),
            .DQ3      ( w_hyper_dq0[3] ),
            .DQ2      ( w_hyper_dq0[2] ),
            .DQ1      ( w_hyper_dq0[1] ),
            .DQ0      ( w_hyper_dq0[0] ),
            .RWDS     ( w_hyper_rwds0  ),
            .CSNeg    ( w_hyper_csn1   ),
            .CK       ( w_hyper_ck     ),
            .CKNeg    ( w_hyper_ckn    ),
            .RESETNeg ( w_hyper_reset  )
         );
         s26ks512s #(
            .TimingModel   ( "S26KS512SDPBHI000"),
            .mem_file_name ( "./vectors/hyper_stim.slm" )
         ) hyperflash_model (
            .DQ7      ( w_hyper_dq0[7] ),
            .DQ6      ( w_hyper_dq0[6] ),
            .DQ5      ( w_hyper_dq0[5] ),
            .DQ4      ( w_hyper_dq0[4] ),
            .DQ3      ( w_hyper_dq0[3] ),
            .DQ2      ( w_hyper_dq0[2] ),
            .DQ1      ( w_hyper_dq0[1] ),
            .DQ0      ( w_hyper_dq0[0] ),
            .RWDS     ( w_hyper_rwds0  ),
            .CSNeg    ( w_hyper_csn0   ),
            .CK       ( w_hyper_ck     ),
            .CKNeg    ( w_hyper_ckn    ),
            .RESETNeg ( w_hyper_reset  )
         );
      end
   endgenerate

   uart_bus #(.BAUD_RATE(115200), .PARITY_EN(0)) i_uart_bus (.rx(w_cva6_uart_tx), .tx(w_cva6_uart_rx), .rx_en(1'b1));

`ifdef SPIKE_TANDEM
    spike #(
        .Size ( NUM_WORDS * 8 )
    ) i_spike (
        .clk_i,
        .rst_ni,
        .clint_tick_i   ( rtc_i                               ),
        .commit_instr_i ( dut.i_ariane.commit_instr_id_commit ),
        .commit_ack_i   ( dut.i_ariane.commit_ack             ),
        .exception_i    ( dut.i_ariane.ex_commit              ),
        .waddr_i        ( dut.i_ariane.waddr_commit_id        ),
        .wdata_i        ( dut.i_ariane.wdata_commit_id        ),
        .priv_lvl_i     ( dut.i_ariane.priv_lvl               )
    );
    initial begin
        $display("Running binary in tandem mode");
    end
`endif

    // Clock process
    initial begin
        clk_i = 1'b0;
        rst_ni = 1'b0;
        repeat(8)
            #(CLOCK_PERIOD/2) clk_i = ~clk_i;
        rst_ni = 1'b1;
        forever begin
            #(CLOCK_PERIOD/2) clk_i = 1'b1;
            #(CLOCK_PERIOD/2) clk_i = 1'b0;

            //if (cycles > max_cycles)
            //    $fatal(1, "Simulation reached maximum cycle count of %d", max_cycles);

            cycles++;
        end
    end

    initial begin
        forever begin
            rtc_i = 1'b0;
            #(RTC_CLOCK_PERIOD/2) rtc_i = 1'b1;
            #(RTC_CLOCK_PERIOD/2) rtc_i = 1'b0;
        end
    end

    initial begin
        forever begin

            wait (exit_o[0]);

            if ((exit_o >> 1)) begin
                `uvm_error( "Core Test",  $sformatf("*** FAILED *** (tohost = %0d)", (exit_o >> 1)))
            end else begin
                `uvm_info( "Core Test",  $sformatf("*** SUCCESS *** (tohost = %0d)", (exit_o >> 1)), UVM_LOW)
            end

            $finish();
        end
    end

    // for faster simulation we can directly preload the ELF
    // Note that we are loosing the capabilities to use risc-fesvr though
    // TODO : preload the ELF on the hyperram instead of the legacy DRAM
    initial begin
        automatic logic [7:0][7:0] mem_row;
        longint address, len;
        byte buffer[];
        void'(uvcl.get_arg_value("+PRELOAD=", binary));

        if (binary != "") begin
            `uvm_info( "Core Test", $sformatf("Preloading ELF: %s", binary), UVM_LOW)

            void'(read_elf(binary));
            // wait with preloading, otherwise randomization will overwrite the existing value
            wait(rst_ni);

           
            // while there are more sections to process
            while (get_section(address, len)) begin
                automatic int num_words = (len+7)/8;
                `uvm_info( "Core Test", $sformatf("Loading Address: %x, Length: %x", address, len),
UVM_LOW)
                buffer = new [num_words*8];
                void'(read_section(address, buffer));
                // preload memories
                // 64-bit
                for (int i = 0; i < num_words; i++) begin
                    mem_row = '0;
                    for (int j = 0; j < 8; j++) begin
                        mem_row[j] = buffer[i*8 + j];
                    end
                end
            end
        end
    end
endmodule // ariane_tb

