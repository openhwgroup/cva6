// Copyright 2021 Thales DIS design services SAS
//
// Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.0
// You may obtain a copy of the License at https://solderpad.org/licenses/
//
// Original Author: Jean-Roch COULON (jean-roch.coulon@thalesgroup.com)


package cva6_config_pkg;

    localparam CVA6ConfigXlen = 32;
    localparam CVA6ConfigFpuEn = 1;
    localparam CVA6ConfigCvxifEn = 0;
    localparam CVA6ConfigCExtEn = 1;

endpackage
