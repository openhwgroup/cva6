// Copyright 2023 Thales
// Copyright 2023 OpenHW Group
//
// Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.0
// You may obtain a copy of the License at https://solderpad.org/licenses/
//
// Original Author: Ayoub JALALI (ayoub.jalali@external.thalesgroup.com)
// ------------------------------------------------------------------------------ //

`DEFINE_ZICOND_INSTR(CZERO_EQZ,        R_FORMAT,  ARITHMETIC, RV32X)
`DEFINE_ZICOND_INSTR(CZERO_NEZ,        R_FORMAT,  ARITHMETIC, RV32X)
