package ariane_pkg;


endpackage