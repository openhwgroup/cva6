// COPYRIGHT HEADER


`ifndef __UVML_SB_MACROS_SV__
`define __UVML_SB_MACROS_SV__





`endif // __UVML_SB_MACROS_SV__
