/*
 * Copyright 2019 Google LLC
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *      http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

//-----------------------------------------------------------------------------
// Processor feature configuration
//-----------------------------------------------------------------------------
// XLEN
parameter int XLEN = 32;

// Parameter for SATP mode, set to BARE if address translation is not supported
parameter satp_mode_t SATP_MODE = BARE;

// Supported Privileged mode
privileged_mode_t supported_privileged_mode[] = {MACHINE_MODE};

// Unsupported instructions
riscv_instr_name_t unsupported_instr[];

// ISA supported by the processor
riscv_instr_group_t supported_isa[$] = {RV32I,
                                        RV32M,
                                        RV32C,
                                        RV32ZBA,
                                        RV32ZBB,
                                        RV32ZBC,
                                        RV32ZBS,
                                        RV32X};

// Interrupt mode support
mtvec_mode_t supported_interrupt_mode[$] = {DIRECT, VECTORED};

// The number of interrupt vectors to be generated, only used if VECTORED interrupt mode is
// supported
int max_interrupt_vector_num = 16;

// Physical memory protection support
bit support_pmp = 0;

// Enhanced physical memory protection support
bit support_epmp = 0;

// Debug mode support
bit support_debug_mode = 0;

// Support delegate trap to user mode
bit support_umode_trap = 0;

// Support sfence.vma instruction
bit support_sfence = 0;

// Support unaligned load/store
bit support_unaligned_load_store = 1'b1;

// GPR setting
parameter int NUM_FLOAT_GPR = 32;
parameter int NUM_GPR = 32;
parameter int NUM_VEC_GPR = 32;

// ----------------------------------------------------------------------------
// Vector extension configuration
// ----------------------------------------------------------------------------

// Parameter for vector extension
parameter int VECTOR_EXTENSION_ENABLE = 0;

parameter int VLEN = 512;

// Maximum size of a single vector element
parameter int ELEN = 32;

// Minimum size of a sub-element, which must be at most 8-bits.
parameter int SELEN = 8;

// Maximum size of a single vector element (encoded in vsew format)
parameter int VELEN = int'($ln(ELEN)/$ln(2)) - 3;

// Maximum LMUL supported by the core
parameter int MAX_LMUL = 8;

// ----------------------------------------------------------------------------
// Multi-harts configuration
// ----------------------------------------------------------------------------

// Number of harts
parameter int NUM_HARTS = 1;

// ----------------------------------------------------------------------------
// Privileged CSR implementation
// ----------------------------------------------------------------------------

// Implemented privileged CSR list
`ifdef DSIM
privileged_reg_t implemented_csr[] = {
`else
const privileged_reg_t implemented_csr[] = {
`endif
    // Machine mode mode CSR
    MVENDORID,        // Vendor ID
    MSTATUS,          // Machine status
    MSTATUSH,         // Additional machine status register, RV32 only
    MISA,             // ISA and extensions
    MIE,              // Machine interrupt-enable register
    MTVEC,            // Machine trap-handler base address
    MSCRATCH,         // Scratch register for machine trap handlers
    MEPC,             // Machine exception program counter
    MCAUSE,           // Machine trap cause
    MTVAL,            // Machine bad address or instruction
    MIP,              // Machine interrupt pending
    MCYCLE,           // Machine cycle counter
    MCYCLEH,          // Upper 32 bits of MCYCLE, RV32I only
    MINSTRETH,        // Upper 32 bits of MINSTRET, RV32I only
    MINSTRET,         // Machine instructions-retired counter
    // Machine Memory Protection
    PMPCFG0,          // Physical memory protection configuration
    PMPCFG1,          // Physical memory protection configuration, RV32 only
    PMPCFG2,          // Physical memory protection configuration
    PMPCFG3,          // Physical memory protection configuration, RV32 only
    PMPADDR0,         // Physical memory protection address register
    PMPADDR1,         // Physical memory protection address register
    PMPADDR2,         // Physical memory protection address register
    PMPADDR3,         // Physical memory protection address register
    PMPADDR4,         // Physical memory protection address register
    PMPADDR5,         // Physical memory protection address register
    PMPADDR6,         // Physical memory protection address register
    PMPADDR7,         // Physical memory protection address register
    PMPADDR8,         // Physical memory protection address register
    PMPADDR9,         // Physical memory protection address register
    PMPADDR10,        // Physical memory protection address register
    PMPADDR11,        // Physical memory protection address register
    PMPADDR12,        // Physical memory protection address register
    PMPADDR13,        // Physical memory protection address register
    PMPADDR14,        // Physical memory protection address register
    PMPADDR15,        // Physical memory protection address register
    // Unprivileged Counter/Timers
    CYCLE,            // Cycle counter for RDCYCLE instruction
    INSTRET,          // Instructions-retired counter for RDINSTRET instruction
    CYCLEH,           // Upper 32 bits of CYCLE, RV32I only
    INSTRETH        // Upper 32 bits of INSTRET, RV32I only
};

// Implementation-specific custom CSRs
bit [11:0] custom_csr[] = {
};

// ----------------------------------------------------------------------------
// Supported interrupt/exception setting, used for functional coverage
// ----------------------------------------------------------------------------

`ifdef DSIM
interrupt_cause_t implemented_interrupt[] = {
`else
const interrupt_cause_t implemented_interrupt[] = {
`endif
    M_SOFTWARE_INTR,
    M_TIMER_INTR,
    M_EXTERNAL_INTR
};

`ifdef DSIM
exception_cause_t implemented_exception[] = {
`else
const exception_cause_t implemented_exception[] = {
`endif
    INSTRUCTION_ADDRESS_MISALIGNED,
    INSTRUCTION_ACCESS_FAULT,
    ILLEGAL_INSTRUCTION,
    BREAKPOINT,
    LOAD_ADDRESS_MISALIGNED,
    LOAD_ACCESS_FAULT,
    STORE_AMO_ADDRESS_MISALIGNED,
    STORE_AMO_ACCESS_FAULT,
    ECALL_MMODE,
    INSTRUCTION_PAGE_FAULT,
    LOAD_PAGE_FAULT,
    STORE_AMO_PAGE_FAULT
};
