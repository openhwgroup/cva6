module scatter_gather(
    input logic    clk,    // Clock
    input logic    aresetn  // Asynchronous reset active low
);

   logic                          dma_req;
   logic                          dma_gnt;
   logic                          dma_rvalid;
   logic                          dma_introut;
   logic [31:0]                   dma_addr;
   logic                          dma_we;
   logic [3:0]                    dma_be;
   logic [31:0]                   dma_rdata;
   logic [31:0]                   dma_wdata;
   logic [31:0]                   dma_tvect;

    AXI_BUS #(
              .AXI_ADDR_WIDTH ( 32 ),
              .AXI_DATA_WIDTH ( 32 ),
              .AXI_ID_WIDTH   ( 4  ),
              .AXI_USER_WIDTH ( 2  )
    ) ctrl_if();
  
core2axi dma_if(
.clk_i(clk),
.rst_ni(aresetn),
.data_req_i(dma_req),
.data_gnt_o(dma_gnt),
.data_rvalid_o(dma_rvalid),
.data_addr_i(dma_addr),
.data_we_i(dma_we),
.data_be_i(dma_be),
.data_rdata_o(dma_rdata),
.data_wdata_i(dma_wdata),

    // ---------------------------------------------------------
    // AXI TARG Port Declarations ------------------------------
    // ---------------------------------------------------------
    //AXI write address bus -------------- // USED// -----------
.aw_id_o(ctrl_if.aw_id),
.aw_addr_o(ctrl_if.aw_addr),
.aw_len_o(ctrl_if.aw_len),
.aw_size_o(ctrl_if.aw_size),
.aw_burst_o(ctrl_if.aw_burst),
.aw_lock_o(ctrl_if.aw_lock),
.aw_cache_o(ctrl_if.aw_cache),
.aw_prot_o(ctrl_if.aw_prot),
.aw_region_o(ctrl_if.aw_region),
.aw_user_o(ctrl_if.aw_user),
.aw_qos_o(ctrl_if.aw_qos),
.aw_valid_o(ctrl_if.aw_valid),
.aw_ready_i(ctrl_if.aw_ready),
    // ---------------------------------------------------------

    //AXI write data bus -------------- // USED// --------------
.w_data_o(ctrl_if.w_data),
.w_strb_o(ctrl_if.w_strb),
.w_last_o(ctrl_if.w_last),
.w_user_o(ctrl_if.w_user),
.w_valid_o(ctrl_if.w_valid),
.w_ready_i(ctrl_if.w_ready),
    // ---------------------------------------------------------

    //AXI write response bus -------------- // USED// ----------
.b_id_i(ctrl_if.b_id),
.b_resp_i(ctrl_if.b_resp),
.b_valid_i(ctrl_if.b_valid),
.b_user_i(ctrl_if.b_user),
.b_ready_o(ctrl_if.b_ready),
    // ---------------------------------------------------------

    //AXI read address bus -------------------------------------
.ar_id_o(ctrl_if.ar_id),
.ar_addr_o(ctrl_if.ar_addr),
.ar_len_o(ctrl_if.ar_len),
.ar_size_o(ctrl_if.ar_size),
.ar_burst_o(ctrl_if.ar_burst),
.ar_lock_o(ctrl_if.ar_lock),
.ar_cache_o(ctrl_if.ar_cache),
.ar_prot_o(ctrl_if.ar_prot),
.ar_region_o(ctrl_if.ar_region),
.ar_user_o(ctrl_if.ar_user),
.ar_qos_o(ctrl_if.ar_qos),
.ar_valid_o(ctrl_if.ar_valid),
.ar_ready_i(ctrl_if.ar_ready),
    // ---------------------------------------------------------

    //AXI read data bus ----------------------------------------
.r_id_i(ctrl_if.r_id),
.r_data_i(ctrl_if.r_data),
.r_resp_i(ctrl_if.r_resp),
.r_last_i(ctrl_if.r_last),
.r_user_i(ctrl_if.r_user),
.r_valid_i(ctrl_if.r_valid),
.r_ready_o(ctrl_if.r_ready)
);

PUMP_AXI4_TO_AXI4 DUT (
	.ARESETn(aresetn),
	.C_CLK(clk),
	.C_ARID(ctrl_if.ar_id),
	.C_ARADDR(ctrl_if.ar_addr),
	.C_ARLEN(ctrl_if.ar_len),
	.C_ARSIZE(ctrl_if.ar_size),
	.C_ARBURST(ctrl_if.ar_burst),
	.C_ARVALID(ctrl_if.ar_valid),
	.C_ARREADY(ctrl_if.ar_ready),
	.C_RID(ctrl_if.r_id),
	.C_RDATA(ctrl_if.r_data),
	.C_RRESP(ctrl_if.r_resp),
	.C_RLAST(ctrl_if.r_last),
	.C_RVALID(ctrl_if.r_valid),
	.C_RREADY(ctrl_if.r_ready),
	.C_AWID(ctrl_if.aw_id),
	.C_AWADDR(ctrl_if.aw_addr),
	.C_AWLEN(ctrl_if.aw_len),
	.C_AWSIZE(ctrl_if.aw_size),
	.C_AWBURST(ctrl_if.aw_burst),
	.C_AWVALID(ctrl_if.aw_valid),
	.C_AWREADY(ctrl_if.aw_ready),
	.C_WDATA(ctrl_if.w_data),
	.C_WSTRB(ctrl_if.w_strb),
	.C_WLAST(ctrl_if.w_last),
	.C_WVALID(ctrl_if.w_valid),
	.C_WREADY(ctrl_if.w_ready),
	.C_BID(ctrl_if.b_id),
	.C_BRESP(ctrl_if.b_resp),
	.C_BVALID(ctrl_if.b_valid),
	.C_BREADY(ctrl_if.b_ready),
	.M_CLK(clk),
	.M_ARID(dbg_master.ar_id),
	.M_ARADDR(dbg_master.ar_addr),
	.M_ARLEN(dbg_master.ar_len),
	.M_ARSIZE(dbg_master.ar_size),
	.M_ARBURST(dbg_master.ar_burst),
	.M_ARLOCK(dbg_master.ar_lock),
	.M_ARCACHE(dbg_master.ar_cache),
	.M_ARPROT(dbg_master.ar_prot),
	.M_ARQOS(dbg_master.ar_qos),
	.M_ARREGION(dbg_master.ar_region),
	.M_ARUSER(dbg_master.ar_user),
	.M_ARVALID(dbg_master.ar_valid),
	.M_ARREADY(dbg_master.ar_ready),
	.M_RID(dbg_master.r_id),
	.M_RDATA(dbg_master.r_data),
	.M_RRESP(dbg_master.r_resp),
	.M_RLAST(dbg_master.r_last),
	.M_RVALID(dbg_master.r_valid),
	.M_RREADY(dbg_master.r_ready),
	.M_AWID(dbg_master.aw_id),
	.M_AWADDR(dbg_master.aw_addr),
	.M_AWLEN(dbg_master.aw_len),
	.M_AWSIZE(dbg_master.aw_size),
	.M_AWBURST(dbg_master.aw_burst),
	.M_AWLOCK(dbg_master.aw_lock),
	.M_AWCACHE(dbg_master.aw_cache),
	.M_AWPROT(dbg_master.aw_prot),
	.M_AWQOS(dbg_master.aw_qos),
	.M_AWREGION(dbg_master.aw_region),
	.M_AWUSER(dbg_master.aw_user),
	.M_AWVALID(dbg_master.aw_valid),
	.M_AWREADY(dbg_master.aw_ready),
	.M_WDATA(dbg_master.w_data),
	.M_WSTRB(dbg_master.w_strb),
	.M_WLAST(dbg_master.w_last),
	.M_WVALID(dbg_master.w_valid),
	.M_WREADY(dbg_master.w_ready),
	.M_BID(dbg_master.b_id),
	.M_BRESP(dbg_master.b_resp),
	.M_BVALID(dbg_master.b_valid),
	.M_BREADY(dbg_master.b_ready),
	.I_CLK(clk),
	.I_ARID(input_if.ar_id),
	.I_ARADDR(input_if.ar_addr),
	.I_ARLEN(input_if.ar_len),
	.I_ARSIZE(input_if.ar_size),
	.I_ARBURST(input_if.ar_burst),
	.I_ARLOCK(input_if.ar_lock),
	.I_ARCACHE(input_if.ar_cache),
	.I_ARPROT(input_if.ar_prot),
	.I_ARQOS(input_if.ar_qos),
	.I_ARREGION(input_if.ar_region),
	.I_ARUSER(input_if.ar_user),
	.I_ARVALID(input_if.ar_valid),
	.I_ARREADY(input_if.ar_ready),
	.I_RID(input_if.r_id),
	.I_RDATA(input_if.r_data),
	.I_RRESP(input_if.r_resp),
	.I_RLAST(input_if.r_last),
	.I_RVALID(input_if.r_valid),
	.I_RREADY(input_if.r_ready),
	.I_AWID(input_if.aw_id),
	.I_AWADDR(input_if.aw_addr),
	.I_AWLEN(input_if.aw_len),
	.I_AWSIZE(input_if.aw_size),
	.I_AWBURST(input_if.aw_burst),
	.I_AWLOCK(input_if.aw_lock),
	.I_AWCACHE(input_if.aw_cache),
	.I_AWPROT(input_if.aw_prot),
	.I_AWQOS(input_if.aw_qos),
	.I_AWREGION(input_if.aw_region),
	.I_AWUSER(input_if.aw_user),
	.I_AWVALID(input_if.aw_valid),
	.I_AWREADY(input_if.aw_ready),
	.I_WDATA(input_if.w_data),
	.I_WSTRB(input_if.w_strb),
	.I_WLAST(input_if.w_last),
	.I_WVALID(input_if.w_valid),
	.I_WREADY(input_if.w_ready),
	.I_BID(input_if.b_id),
	.I_BRESP(input_if.b_resp),
	.I_BVALID(input_if.b_valid),
	.I_BREADY(input_if.b_ready),
	.O_CLK(clk),
	.O_ARID(output_if.ar_id),
	.O_ARADDR(output_if.ar_addr),
	.O_ARLEN(output_if.ar_len),
	.O_ARSIZE(output_if.ar_size),
	.O_ARBURST(output_if.ar_burst),
	.O_ARLOCK(output_if.ar_lock),
	.O_ARCACHE(output_if.ar_cache),
	.O_ARPROT(output_if.ar_prot),
	.O_ARQOS(output_if.ar_qos),
	.O_ARREGION(output_if.ar_region),
	.O_ARUSER(output_if.ar_user),
	.O_ARVALID(output_if.ar_valid),
	.O_ARREADY(output_if.ar_ready),
	.O_RID(output_if.r_id),
	.O_RDATA(output_if.r_data),
	.O_RRESP(output_if.r_resp),
	.O_RLAST(output_if.r_last),
	.O_RVALID(output_if.r_valid),
	.O_RREADY(output_if.r_ready),
	.O_AWID(output_if.aw_id),
	.O_AWADDR(output_if.aw_addr),
	.O_AWLEN(output_if.aw_len),
	.O_AWSIZE(output_if.aw_size),
	.O_AWBURST(output_if.aw_burst),
	.O_AWLOCK(output_if.aw_lock),
	.O_AWCACHE(output_if.aw_cache),
	.O_AWPROT(output_if.aw_prot),
	.O_AWQOS(output_if.aw_qos),
	.O_AWREGION(output_if.aw_region),
	.O_AWUSER(output_if.aw_user),
	.O_AWVALID(output_if.aw_valid),
	.O_AWREADY(output_if.aw_ready),
	.O_WDATA(output_if.w_data),
	.O_WSTRB(output_if.w_strb),
	.O_WLAST(output_if.w_last),
	.O_WVALID(output_if.w_valid),
	.O_WREADY(output_if.w_ready),
	.O_BID(output_if.b_id),
	.O_BRESP(output_if.b_resp),
	.O_BVALID(output_if.b_valid),
	.O_BREADY(output_if.b_ready),
	.I_IRQ(i_irq),
	.O_IRQ(o_irq)
);
 
endmodule
