/*
 * Copyright 2018 Google LLC
 * Copyright 2020 OpenHW Group
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *      http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

//-----------------------------------------------------------------------------
// Copy/Modify version of riscv-dv/tests/riscv_instr_gen_tb_top.sv to add the
// corev specific tests.
//-----------------------------------------------------------------------------
module cv32e40p_instr_gen_tb_top;

  import uvm_pkg::*;
  import riscv_instr_test_pkg::*;
  import corev_instr_test_pkg::*;
  import cv32e40p_instr_test_pkg::*;

  initial begin
    run_test();
  end

endmodule : cv32e40p_instr_gen_tb_top
