package eth_tb_pkg;

    `include "sequence_item.svh"
    `include "driver.svh"

endpackage