`ifndef __UVMA_CVA6PKG_UTILS_PKG_SV__
`define __UVMA_CVA6PKG_UTILS_PKG_SV__

package uvma_cva6pkg_utils_pkg;

    import ariane_pkg::*;
    import cva6_config_pkg::*;
    import uvma_core_cntrl_pkg::*;
   `include "uvma_cva6pkg_utils.sv"

endpackage : uvma_cva6pkg_utils_pkg

`endif
