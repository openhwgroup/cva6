/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 942;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h0a0d2165_6e6f6420,
        64'h00000000_00206567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f63,
        64'h00000000_00000009,
        64'h3a656d61_6e090a0d,
        64'h00093a73_65747562,
        64'h69727474_61090a0d,
        64'h00000009_3a61626c,
        64'h20747361_6c090a0d,
        64'h0000093a_61626c20,
        64'h74737269_66090a0d,
        64'h00000000_00000000,
        64'h09202020_20203a64,
        64'h69756720_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_00000000,
        64'h093a6469_75672065,
        64'h70797420_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20747067,
        64'h00000009_20203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20657a69_73090a0d,
        64'h00000009_3a736569,
        64'h72746e65_206e6f69,
        64'h74697472_61702072,
        64'h65626d75_6e090a0d,
        64'h00000009_2020203a,
        64'h61626c20_73656972,
        64'h746e6520_6e6f6974,
        64'h69747261_70090a0d,
        64'h00093a61_646c2070,
        64'h756b6361_62090a0d,
        64'h00000000_00000000,
        64'h093a6162_6c20746e,
        64'h65727275_63090a0d,
        64'h00000009_3a646576,
        64'h72657365_72090a0d,
        64'h00093a72_65646165,
        64'h685f6372_63090a0d,
        64'h00000000_00000909,
        64'h3a657a69_73090a0d,
        64'h00000009_3a6e6f69,
        64'h73697665_72090a0d,
        64'h0000093a_65727574,
        64'h616e6769_73090a0d,
        64'h00000000_003a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20747067,
        64'h0000203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_63206473,
        64'h00000000_0000000a,
        64'h0d216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_0000000a,
        64'h0d216465_7a696c61,
        64'h6974696e_69206473,
        64'h00000000_0a0d676e,
        64'h69746978_65202e2e,
        64'h2e647320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f63,
        64'h00000000_0000002e,
        64'h0000000a_0d202e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e69,
        64'h00000031_34646d63,
        64'h00000035_35646d63,
        64'h00000000_30646d63,
        64'h00000020_3a206573,
        64'h6e6f7073_65720920,
        64'h00000000_0020646e,
        64'h616d6d6f_63204453,
        64'h00000000_203f3f79,
        64'h74706d65_20746f6e,
        64'h206f6669_66207872,
        64'h00000000_00000a0d,
        64'h2164657a_696c6169,
        64'h74696e69_20495053,
        64'h00000000_00007830,
        64'h203a7375_74617473,
        64'h00000000_00000a0d,
        64'h49505320_74696e69,
        64'h00000a0d_21646c72,
        64'h6f57206f_6c6c6548,
        64'h00000032_2d746c75,
        64'h61666564_2d697274,
        64'h2c786e6c_7800746c,
        64'h75616665_642d6972,
        64'h742c786e_6c78006c,
        64'h6175642d_73692c78,
        64'h6e6c7800_746e6573,
        64'h6572702d_74707572,
        64'h7265746e_692c786e,
        64'h6c780068_74646977,
        64'h2d326f69_70672c78,
        64'h6e6c7800_68746469,
        64'h772d6f69_70672c78,
        64'h6e6c7800_322d746c,
        64'h75616665_642d7475,
        64'h6f642c78_6e6c7800,
        64'h746c7561_6665642d,
        64'h74756f64_2c786e6c,
        64'h7800322d_73747570,
        64'h6e692d6c_6c612c78,
        64'h6e6c7800_73747570,
        64'h6e692d6c_6c612c78,
        64'h6e6c7800_72656c6c,
        64'h6f72746e_6f632d6f,
        64'h69706700_736c6c65,
        64'h632d6f69_70672300,
        64'h6f69646d_2d736168,
        64'h2c786e6c_78006c61,
        64'h6e726574_6e692d65,
        64'h73752c78_6e6c7800,
        64'h676e6f70_2d676e69,
        64'h702d7874_2c786e6c,
        64'h78006874_6469772d,
        64'h64692d69_78612d73,
        64'h2c786e6c_7800676e,
        64'h6f702d67_6e69702d,
        64'h78722c78_6e6c7800,
        64'h65636e61_74736e69,
        64'h2c786e6c_78006f69,
        64'h646d2d65_64756c63,
        64'h6e692c78_6e6c7800,
        64'h6b636162_706f6f6c,
        64'h2d6c616e_7265746e,
        64'h692d6564_756c636e,
        64'h692c786e_6c780073,
        64'h72656666_75622d6c,
        64'h61626f6c_672d6564,
        64'h756c636e_692c786e,
        64'h6c780078_656c7075,
        64'h642c786e_6c780065,
        64'h6c646e61_682d7968,
        64'h70007373_65726464,
        64'h612d6361_6d2d6c61,
        64'h636f6c00_70772d65,
        64'h6c626173_69640073,
        64'h65676e61_722d6567,
        64'h61746c6f_76007963,
        64'h6e657571_6572662d,
        64'h78616d2d_69707300,
        64'h6f697461_722d6b63,
        64'h732c786e_6c780073,
        64'h7469622d_72656673,
        64'h6e617274_2d6d756e,
        64'h2c786e6c_78007374,
        64'h69622d73_732d6d75,
        64'h6e2c786e_6c780074,
        64'h73697865_2d6f6669,
        64'h662c786e_6c780079,
        64'h6c696d61_662c786e,
        64'h6c780068_74646977,
        64'h2d6f692d_67657200,
        64'h74666968_732d6765,
        64'h72007374_70757272,
        64'h65746e69_00746e65,
        64'h7261702d_74707572,
        64'h7265746e_69006465,
        64'h6570732d_746e6572,
        64'h72756300_7665646e,
        64'h2c766373_69720079,
        64'h7469726f_6972702d,
        64'h78616d2c_76637369,
        64'h72007365_6d616e2d,
        64'h67657200_6465646e,
        64'h65747865_2d737470,
        64'h75727265_746e6900,
        64'h7365676e_61720064,
        64'h65646e65_70737573,
        64'h2d657461_74732d6e,
        64'h69617465_72007265,
        64'h67676972_742d746c,
        64'h75616665_642c7875,
        64'h6e696c00_736f6970,
        64'h6700656c_646e6168,
        64'h702c7875_6e696c00,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_00736c6c,
        64'h65632d74_70757272,
        64'h65746e69_23007469,
        64'h6c70732d_626c7400,
        64'h65707974_2d756d6d,
        64'h00617369_2c766373,
        64'h69720073_75746174,
        64'h73006765_72006570,
        64'h79745f65_63697665,
        64'h64007963_6e657571,
        64'h6572662d_6b636f6c,
        64'h63007963_6e657571,
        64'h6572662d_65736162,
        64'h656d6974_00687461,
        64'h702d7475_6f647473,
        64'h006c6564_6f6d0065,
        64'h6c626974_61706d6f,
        64'h6300736c_6c65632d,
        64'h657a6973_2300736c,
        64'h6c65632d_73736572,
        64'h64646123_09000000,
        64'h02000000_02000000,
        64'h02000000_01000000,
        64'hbb000000_04000000,
        64'h03000000_01000000,
        64'hb5000000_04000000,
        64'h03000000_ffffffff,
        64'h8f030000_04000000,
        64'h03000000_ffffffff,
        64'h7e030000_04000000,
        64'h03000000_01000000,
        64'h71030000_04000000,
        64'h03000000_00000000,
        64'h5a030000_04000000,
        64'h03000000_08000000,
        64'h49030000_04000000,
        64'h03000000_08000000,
        64'h39030000_04000000,
        64'h03000000_00000000,
        64'h25030000_04000000,
        64'h03000000_00000000,
        64'h13030000_04000000,
        64'h03000000_00000000,
        64'h01030000_04000000,
        64'h03000000_00000000,
        64'hf1020000_04000000,
        64'h03000000_00000100,
        64'h00000000_00000040,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'he1020000_00000000,
        64'h03000000_00000000,
        64'h612e3030_2e312d6f,
        64'h6970672d_7370782c,
        64'h786e6c78_1b000000,
        64'h15000000_03000000,
        64'h02000000_d5020000,
        64'h04000000_03000000,
        64'h00000030_30303030,
        64'h30303440_6f697067,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h04000000_bb000000,
        64'h04000000_03000000,
        64'h04000000_b5000000,
        64'h04000000_03000000,
        64'h01000000_67000000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_00000000,
        64'h35313943_2e433130,
        64'h3064692d_7968702d,
        64'h74656e72_65687465,
        64'h1b000000_19000000,
        64'h03000000_00000031,
        64'h406f6964_6d5f305f,
        64'h6574696c_74656e72,
        64'h65687465_5f697861,
        64'h01000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h6f69646d_01000000,
        64'h01000000_c7020000,
        64'h04000000_03000000,
        64'h00000000_b5020000,
        64'h04000000_03000000,
        64'h01000000_a3020000,
        64'h04000000_03000000,
        64'h04000000_8f020000,
        64'h04000000_03000000,
        64'h01000000_7d020000,
        64'h04000000_03000000,
        64'h00657469_6c74656e,
        64'h72656874_655f6978,
        64'h615f786e_6c785f69,
        64'h6f020000_18000000,
        64'h03000000_01000000,
        64'h5d020000_04000000,
        64'h03000000_00000000,
        64'h3e020000_04000000,
        64'h03000000_01000000,
        64'h22020000_04000000,
        64'h03000000_01000000,
        64'h16020000_04000000,
        64'h03000000_00000100,
        64'h00000000_00000030,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h04000000_0b020000,
        64'h04000000_03000000,
        64'h00002201_00350a00,
        64'hf9010000_06000000,
        64'h03000000_00000000,
        64'h03000000_58010000,
        64'h08000000_03000000,
        64'h03000000_47010000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_0000612e,
        64'h30302e31_2d657469,
        64'h6c74656e_72656874,
        64'h652d7370_782c786e,
        64'h6c780030_2e332d65,
        64'h74696c74_656e7265,
        64'h6874652d_6978612c,
        64'h786e6c78_1b000000,
        64'h37000000_03000000,
        64'h00000030_30303030,
        64'h30303340_74656e72,
        64'h65687465_01000000,
        64'h02000000_02000000,
        64'hee010000_00000000,
        64'h03000000_e40c0000,
        64'he40c0000_df010000,
        64'h08000000_03000000,
        64'h20bcbe00_cd010000,
        64'h04000000_03000000,
        64'h00000000_67000000,
        64'h04000000_03000000,
        64'h00000000_746f6c73,
        64'h2d697073_2d636d6d,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h40636d6d_01000000,
        64'h04000000_be010000,
        64'h04000000_03000000,
        64'h08000000_a7010000,
        64'h04000000_03000000,
        64'h01000000_96010000,
        64'h04000000_03000000,
        64'h01000000_86010000,
        64'h04000000_03000000,
        64'h00377865_746e696b,
        64'h7a010000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h02000000_02000000,
        64'h58010000_08000000,
        64'h03000000_03000000,
        64'h47010000_04000000,
        64'h03000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_00612e30,
        64'h302e322d_6970732d,
        64'h7370782c_786e6c78,
        64'h00622e30_302e322d,
        64'h6970732d_7370782c,
        64'h786e6c78_1b000000,
        64'h28000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40697073,
        64'h2d737078_01000000,
        64'h02000000_04000000,
        64'h6d010000_04000000,
        64'h03000000_02000000,
        64'h63010000_04000000,
        64'h03000000_01000000,
        64'h58010000_04000000,
        64'h03000000_03000000,
        64'h47010000_04000000,
        64'h03000000_00c20100,
        64'h39010000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000010,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00303537_3631736e,
        64'h1b000000_08000000,
        64'h03000000_00000030,
        64'h30303030_30303140,
        64'h74726175_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_11010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000000_00000000,
        64'h67000000_10000000,
        64'h03000000_ffff0000,
        64'h02000000_fd000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00003040,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h03000000_bb000000,
        64'h04000000_03000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h03000000_2e010000,
        64'h04000000_03000000,
        64'h07000000_1b010000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h02000000_0b000000,
        64'h02000000_fd000000,
        64'h10000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_11010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_fd000000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hf6000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_02000000,
        64'hdf000000_00000000,
        64'h03000000_00000074,
        64'h61656274_72616568,
        64'hc9000000_0a000000,
        64'h03000000_00000000,
        64'h01000000_01000000,
        64'hc3000000_0c000000,
        64'h03000000_00000064,
        64'h656c2d74_61656274,
        64'h72616568_01000000,
        64'h00000073_64656c2d,
        64'h6f697067_1b000000,
        64'h0a000000_03000000,
        64'h00000000_7364656c,
        64'h01000000_02000000,
        64'h00000008_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_bb000000,
        64'h04000000_03000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00007573_63616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hac0a0000_a2030000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'he40a0000_38000000,
        64'h860e0000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'ha0018402_19c58593,
        64'h00000597_01f41413,
        64'h0010041b_e911d31f,
        64'hf0ef057e_65a14505,
        64'hf16ff0ef_04450513,
        64'h00001517_ef0ff0ef,
        64'he4061141_bbb5f2cf,
        64'hf0ef32a5_05130000,
        64'h1517b3f5_0a450513,
        64'h00001517_fc4ff0ef,
        64'h8526f48f_f0ef1865,
        64'h05130000_1517f54f,
        64'hf0ef17a5_05130000,
        64'h1517c50d_84aac5ff,
        64'hf0ef8552_865a020a,
        64'ha583f70f_f0ef3565,
        64'h05130000_1517f579,
        64'h93e30804_8493f84f,
        64'hf0ef2985_0f450513,
        64'h00001517_ff2c1be3,
        64'h85bff0ef_09050009,
        64'h4503fa0f_f0ef3765,
        64'h05130000_151782ff,
        64'hf0ef7088_fb2ff0ef,
        64'h37850513_00001517,
        64'h841ff0ef_6c88fc4f,
        64'hf0ef37a5_05130000,
        64'h1517853f_f0ef0704,
        64'h8c130284_89136888,
        64'hfdeff0ef_38450513,
        64'h00001517_ff2c1be3,
        64'h8b3ff0ef_09050009,
        64'h45030109_0c13ffcf,
        64'hf0ef3825_05130000,
        64'h1517fe99_1be38d1f,
        64'hf0ef0905_00094503,
        64'hff048913_81bff0ef,
        64'h38050513_00001517,
        64'h8ebff0ef_0ff9f513,
        64'h82fff0ef_37c50513,
        64'h00001517_b5fd1a65,
        64'h05130000_15178c7f,
        64'hf0ef854e_84bff0ef,
        64'h28850513_00001517,
        64'h857ff0ef_27c50513,
        64'h00001517_c50d0804,
        64'h89aa8a8a_d65ff0ef,
        64'h850a4605_71010489,
        64'h2583879f_f0ef1e65,
        64'h05130000_15178c7f,
        64'hf0ef4556_88bff0ef,
        64'h3b850513_00001517,
        64'h8d9ff0ef_454689df,
        64'hf0ef3aa5_05130000,
        64'h151792bf_f0ef6526,
        64'h8afff0ef_39c50513,
        64'h00001517_93dff0ef,
        64'h75028c1f_f0ef39e5,
        64'h05130000_151794ff,
        64'hf0ef6562_8d3ff0ef,
        64'h39850513_00001517,
        64'h921ff0ef_45528e5f,
        64'hf0ef39a5_05130000,
        64'h1517933f_f0ef4542,
        64'h8f7ff0ef_39c50513,
        64'h00001517_945ff0ef,
        64'h4532909f_f0ef39e5,
        64'h05130000_1517957f,
        64'hf0ef4522_91bff0ef,
        64'h3a050513_00001517,
        64'h9a9ff0ef_4b916502,
        64'h92fff0ef_3a450513,
        64'h00001517_93bff0ef,
        64'h39050513_00001517,
        64'hbf6154f9_94bff0ef,
        64'h2b850513_00001517,
        64'h9d9ff0ef_852695df,
        64'hf0ef39a5_05130000,
        64'h1517969f_f0ef38e5,
        64'h05130000_1517c905,
        64'h84aa890a_e75ff0ef,
        64'h850a4585_46057101,
        64'h987ff0ef_39450513,
        64'h00001517_80826161,
        64'h6c026ba2_6b426ae2,
        64'h7a0279a2_794274e2,
        64'h64068526_60a6fb04,
        64'h011354fd_9b3ff0ef,
        64'h39850513_00001517,
        64'hc51de1ff_f0ef8b2e,
        64'h8a2a0880_e062e45e,
        64'hec56f44e_f84afc26,
        64'he486e85a_f052e0a2,
        64'h715dbfe1_54798082,
        64'h61696baa_6b4a6aea,
        64'h7a0a79aa_794a74ea,
        64'h640e60ae_8522c77f,
        64'hf0efc83f_f0ef4531,
        64'h45814605_4401f890,
        64'h46e314fd_a13ff0ef,
        64'h3f050513_00001517,
        64'he7990354_e7b30534,
        64'h12632981_90411442,
        64'h8c49cabf_f0ef9041,
        64'h03051413_89220085,
        64'h151bcbbf_f0effd64,
        64'h1ae30404_0413ff79,
        64'h17e389aa_f0fff0ef,
        64'h0905854e_0007c583,
        64'h012407b3_04000b93,
        64'h4901c63f_f0ef850a,
        64'h04000593_86224981,
        64'h844a2009_0b13ff45,
        64'h1ee3cfbf_f0ef3e80,
        64'h0a930fe0_0a139081,
        64'h1482bff5_d0dff0ef,
        64'hc501d1bf_f0ef4549,
        64'h85a20ff6_76130016,
        64'h66130015_161bf4ff,
        64'hf0ef0ff4_7593f57f,
        64'hf0ef0ff5_f5930084,
        64'h559bf63f_f0ef0ff5,
        64'hf5930104_559bf6ff,
        64'hf0ef4501_0ff5f593,
        64'h0184559b_fee79be3,
        64'h078500c6_802300f1,
        64'h06b30800_0713567d,
        64'h4781842e_892ae55e,
        64'he95aed56_f152f54e,
        64'he58684b2_f94afd26,
        64'he1a27155_80829141,
        64'h15428d3d_8ff90057,
        64'h979b1701_67090107,
        64'hd79b0105_179b4105,
        64'h551b0105_151b8d2d,
        64'h00c59513_8da9893d,
        64'h0045d51b_8da99141,
        64'h15428d5d_05220085,
        64'h579b8082_07f57513,
        64'h8d2d0045_15938d2d,
        64'h8d3d0045_d51b0075,
        64'hd79b8de9_80820141,
        64'h853e6402_60a24781,
        64'hc11157f5_f89ff0ef,
        64'hc51157f9_efbff0ef,
        64'hc91157fd_eb7ff0ef,
        64'hfc6de03f_f0ef347d,
        64'h4429b91f_f0ef5565,
        64'h05130000_1517c89f,
        64'hf0efe022_e4061141,
        64'h80826105_00153513,
        64'h64a26442_60e20004,
        64'h051bfc94_0ce3e37f,
        64'hf0efeb3f_f0ef57e5,
        64'h05130000_151785aa,
        64'h842ae53f_f0ef0290,
        64'h05134000_05b70770,
        64'h0613fbdf_f0ef4485,
        64'he822ec06_e4261101,
        64'h80820141_00153513,
        64'h157d6402_60a20004,
        64'h051bef3f_f0ef5b85,
        64'h051385a2_00001517,
        64'he89ff0ef_842ae97f,
        64'hf0efe022_e4060370,
        64'h05134581_06500613,
        64'h11418082_61056902,
        64'h64a26442_60e20015,
        64'h3513f565_05130004,
        64'h051b0124_986388bd,
        64'h00f91b63_45014785,
        64'hec9ff0ef_ecdff0ef,
        64'h842aed3f_f0ef84aa,
        64'hed9ff0ef_eddff0ef,
        64'hee1ff0ef_892aeeff,
        64'hf0efe04a_e426e822,
        64'hec064521_1aa00593,
        64'h08700613_1101bfcd,
        64'h45018082_61056902,
        64'h64a26442_60e24505,
        64'hf89ff0ef_45856465,
        64'h05130000_1517fe99,
        64'h15e3c00d_f25ff0ef,
        64'h892a347d_f35ff0ef,
        64'h45014581_09500613,
        64'h44857104_0413e04a,
        64'hec06e426_6409e822,
        64'h1101cd1f_f06f6105,
        64'h64050513_00001517,
        64'h60e26442_da7ff0ef,
        64'h852e65a2_cebff0ef,
        64'h68850513_00001517,
        64'hcf7ff0ef_8522cfdf,
        64'hf0efe42e_ec0668e5,
        64'h05130000_1517842a,
        64'he8221101_80826145,
        64'h64e27402_70a2f47d,
        64'h147d0007_d4634187,
        64'hd79b0185_179bfa7f,
        64'hf0efeb5f_f0ef8532,
        64'h06400413_6622ec1f,
        64'hf0ef0ff4_7513ec9f,
        64'hf0ef0ff5_75130084,
        64'h551bed5f_f0ef0ff5,
        64'h75130104_551bee1f,
        64'hf0ef0ff5_75130184,
        64'h551beedf_f0ef0404,
        64'he513febf_f0ef84aa,
        64'h842eec26_f022e432,
        64'hf4067179_f07ff06f,
        64'h0ff00513_8082557d,
        64'hb7e900d7_00230785,
        64'h00f60733_06c82683,
        64'hff798b05_5178bf4d,
        64'hd6b80785_0007c703,
        64'h80824501_d3b84719,
        64'hdbb8577d_200007b7,
        64'h00b6ef63_0007869b,
        64'h20000837_20000537,
        64'hfff58b85_537c2000,
        64'h0737d3b8_200007b7,
        64'h10600713_fff537fd,
        64'h00010320_079304b7,
        64'h616340a7_873b87aa,
        64'h200006b7_dbb85779,
        64'h200007b7_06b7ec63,
        64'h10000793_80826105,
        64'h64a2d3b8_4719dbb8,
        64'h644260e2_0ff47513,
        64'h577d2000_07b7e25f,
        64'hf0ef7925_05130000,
        64'h1517eb3f_f0ef9101,
        64'h15024088_e3bff0ef,
        64'h7b050513_00001517,
        64'he3958b85_240153fc,
        64'h57e0ff65_8b050647,
        64'h849353f8_d3b81060,
        64'h07132000_07b7fff5,
        64'h37fd0001_06400793,
        64'hd7a8dbb8_5779e426,
        64'he822ec06_200007b7,
        64'h1101e81f_f06f6105,
        64'h7e050513_00001517,
        64'h64a260e2_6442d03c,
        64'h4799e99f_f0ef8065,
        64'h05130000_2517f27f,
        64'hf0ef9101_02049513,
        64'h2481eb1f_f0ef7fe5,
        64'h05130000_15175064,
        64'hd03c1660_0793ec5f,
        64'hf0ef8325_05130000,
        64'h2517f53f_f0ef9101,
        64'h02049513_2481eddf,
        64'hf0ef82a5_05130000,
        64'h25175064_d03c1040,
        64'h07932000_0437fff5,
        64'h37fd0001_47a9c3b8,
        64'h47292000_07b7f05f,
        64'hf0efe426_e822ec06,
        64'h84a50513_11010000,
        64'h25178082_41088082,
        64'hc10c8082_610560e2,
        64'hee1ff0ef_00914503,
        64'hee9ff0ef_00814503,
        64'hf55ff0ef_ec06002c,
        64'h11018082_61456942,
        64'h64e27402_70a2fe94,
        64'h10e3f0bf_f0ef0091,
        64'h4503f13f_f0ef3461,
        64'h00814503_f81ff0ef,
        64'h0ff57513_002c0089,
        64'h553354e1_03800413,
        64'h892af406_e84aec26,
        64'hf0227179_80826145,
        64'h694264e2_740270a2,
        64'hfe9410e3_f4dff0ef,
        64'h00914503_f55ff0ef,
        64'h34610081_4503fc3f,
        64'hf0ef0ff5_7513002c,
        64'h0089553b_54e14461,
        64'h892af406_e84aec26,
        64'hf0227179_808200f5,
        64'h80230007_c78300e5,
        64'h80a397aa_81110007,
        64'h4703973e_00f57713,
        64'h98078793_00001797,
        64'hb7f50405_fa5ff0ef,
        64'h80820141_640260a2,
        64'he5090004_4503842a,
        64'he406e022_11418082,
        64'h00e78823_02000713,
        64'h00e78423_fc700713,
        64'h00e78623_470d0007,
        64'h822300e7_8023476d,
        64'h00e78623_f8000713,
        64'h00078223_100007b7,
        64'h808200a7_0023dfe5,
        64'h0207f793_01474783,
        64'h10000737_80820205,
        64'h75130147_c5031000,
        64'h07b78082_00054503,
        64'h808200b5_00238082,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_01f49493,
        64'h0010049b_b8458593,
        64'h00001597_f1402573,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'hfe091ee3_0004a903,
        64'h00092023_00990933,
        64'h00291913_f1402973,
        64'h020004b7_fe090ae3,
        64'h00897913_34402973,
        64'h10500073_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_0124a023,
        64'h00100913_020004b7,
        64'h221000ef_01a11113,
        64'h0210011b_03249663,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
