/*
 *
 * Copyright (c) 2005-2020 Imperas Software Ltd., www.imperas.com
 *
 * The contents of this file are provided under the Software License 
 * Agreement that you accepted before downloading this file.
 *
 * This source forms part of the Software and can be used for educational,
 * training, and demonstration purposes but cannot be used for derivative
 * works except in cases where the derivative works require OVP technology
 * to run. 
 *
 * For open source models released under licenses that you can use for 
 * derivative works, please visit www.OVPworld.org or www.imperas.com
 * for the location of the open source models. 
 *
 */

// Coverage for : RVI,RVIpseudo

// This file is auto generated by Imperas.
// It is an example of SystemVerilog UVM functional coverage.

typedef enum {
    ADD,ADDI,AND,ANDI,AUIPC,BEQ,BEQZ,BGE,BGEU,
    BGEZ,BGTZ,BLEZ,BLT,BLTU,BLTZ,BNE,BNEZ,
    EBREAK,ECALL,ILLEGAL,J,JAL,JALR,JR,LB,
    LBU,LH,LHU,LUI,LW,MV,NEG,NOP,
    NOT,OR,ORI,RET,SB,SEQZ,SGTZ,SH,
    SLL,SLLI,SLT,SLTI,SLTIU,SLTU,SLTZ,SNEZ,
    SRA,SRAI,SRL,SRLI,SUB,SW,XOR,XORI,
    CSRW,
    NOT_YET_INCLUDED
} instr_name_t;

typedef struct {
    string key;
    string val;
} ops_t;

typedef struct {
    string ins_str;
    instr_name_t asm;
    ops_t ops[4];
} ins_t;

class coverage;

    function instr_name_t get_asm_enum(string ins_str);
        case (ins_str)
            "add": return ADD;
            "addi": return ADDI;
            "and": return AND;
            "andi": return ANDI;
            "auipc": return AUIPC;
            "beq": return BEQ;
            "beqz": return BEQZ;
            "bge": return BGE;
            "bgeu": return BGEU;
            "bgez": return BGEZ;
            "bgtz": return BGTZ;
            "blez": return BLEZ;
            "blt": return BLT;
            "bltu": return BLTU;
            "bltz": return BLTZ;
            "bne": return BNE;
            "bnez": return BNEZ;
            "ebreak": return EBREAK;
            "ecall": return ECALL;
            "illegal": return ILLEGAL;
            "j": return J;
            "jal": return JAL;
            "jalr": return JALR;
            "jr": return JR;
            "lb": return LB;
            "lbu": return LBU;
            "lh": return LH;
            "lhu": return LHU;
            "lui": return LUI;
            "lw": return LW;
            "mv": return MV;
            "neg": return NEG;
            "nop": return NOP;
            "not": return NOT;
            "or": return OR;
            "ori": return ORI;
            "ret": return RET;
            "sb": return SB;
            "seqz": return SEQZ;
            "sgtz": return SGTZ;
            "sh": return SH;
            "sll": return SLL;
            "slli": return SLLI;
            "slt": return SLT;
            "slti": return SLTI;
            "sltiu": return SLTIU;
            "sltu": return SLTU;
            "sltz": return SLTZ;
            "snez": return SNEZ;
            "sra": return SRA;
            "srai": return SRAI;
            "srl": return SRL;
            "srli": return SRLI;
            "sub": return SUB;
            "sw": return SW;
            "xor": return XOR;
            "xori": return XORI;
            "csrw": return CSRW;
            default: begin
                $display("ERROR: get_asm_enum(%0s) not found in enum list", ins_str);
                //$finish(-1);
            end
        endcase
    endfunction

    covergroup ins_cg with function sample(string ins_str);
        option.per_instance = 1;
        cp_asm : coverpoint get_asm_enum(ins_str);
    endgroup

    function new();
        ins_cg = new();
    endfunction

    function void sample(input string decode);
        string ins_str, op[4], key, val;
        int num = $sscanf (decode, "%s %s %s %s %s", ins_str, op[0], op[1], op[2], op[3]);
        ins_cg.sample(ins_str);
    endfunction

endclass
