// COPYRIGHT HEADER


`ifndef __UVML_HRTBT_CONSTANTS_SV__
`define __UVML_HRTBT_CONSTANTS_SV__





`endif // __UVML_HRTBT_CONSTANTS_SV__
