module hpdcache_priv_adapter
  import ariane_pkg::*;
  #(parameter config_pkg::cva6_cfg_t CVA6Cfg = config_pkg::cva6_cfg_empty,
    parameter type icache_areq_t = logic,
    parameter type icache_arsp_t = logic,
    parameter type icache_dreq_t = logic,
    parameter type icache_drsp_t = logic,
    parameter type icache_req_t = logic,
    parameter type icache_rtrn_t = logic,
    parameter type dcache_req_i_t = logic,
    parameter type dcache_req_o_t = logic,
    parameter int NumPorts = 4,
    parameter int NrHwPrefetchers = 4,
    parameter type axi_ar_chan_t = logic,
    parameter type axi_aw_chan_t = logic,
    parameter type axi_w_chan_t = logic,
    parameter type axi_b_chan_t = logic,
    parameter type axi_r_chan_t = logic,
    parameter type noc_req_t = logic,
    parameter type noc_resp_t = logic,
    parameter type cmo_req_t = logic,
    parameter type cmo_rsp_t = logic)
   (
    input logic clk_i,
    input logic rst_ni,
    input riscv::priv_lvl_t priv_lvl_i,
    output noc_req_t  noc_req_o,
    input  noc_resp_t noc_resp_i,
    input logic icache_en_i,
    input logic icache_flush_i,
    output logic icache_miss_o,
    input icache_areq_t icache_areq_i,
    output icache_arsp_t icache_areq_o,
    input icache_dreq_t icache_dreq_i,
    output icache_drsp_t icache_dreq_o,
    input  logic dcache_enable_i,
    input  logic dcache_flush_i,
    output logic dcache_flush_ack_o,
    output logic dcache_miss_o,
    input  ariane_pkg::amo_req_t dcache_amo_req_i,
    output ariane_pkg::amo_resp_t dcache_amo_resp_o,
    input  cmo_req_t dcache_cmo_req_i,
    output cmo_rsp_t dcache_cmo_resp_o,
    input  dcache_req_i_t [NumPorts-1:0] dcache_req_ports_i,
    output dcache_req_o_t [NumPorts-1:0] dcache_req_ports_o,
    output logic wbuffer_empty_o,
    output logic wbuffer_not_ni_o,
    input  logic [NrHwPrefetchers-1:0]       hwpf_base_set_i,
    input  logic [NrHwPrefetchers-1:0][63:0] hwpf_base_i,
    output logic [NrHwPrefetchers-1:0][63:0] hwpf_base_o,
    input  logic [NrHwPrefetchers-1:0]       hwpf_param_set_i,
    input  logic [NrHwPrefetchers-1:0][63:0] hwpf_param_i,
    output logic [NrHwPrefetchers-1:0][63:0] hwpf_param_o,
    input  logic [NrHwPrefetchers-1:0]       hwpf_throttle_set_i,
    input  logic [NrHwPrefetchers-1:0][63:0] hwpf_throttle_i,
    output logic [NrHwPrefetchers-1:0][63:0] hwpf_throttle_o,
    output logic [63:0] hwpf_status_o
   );
   cva6_hpdcache_subsystem #(
     .CVA6Cfg(CVA6Cfg),
     .icache_areq_t(icache_areq_t),
     .icache_arsp_t(icache_arsp_t),
     .icache_dreq_t(icache_dreq_t),
     .icache_drsp_t(icache_drsp_t),
     .icache_req_t(icache_req_t),
     .icache_rtrn_t(icache_rtrn_t),
     .dcache_req_i_t(dcache_req_i_t),
     .dcache_req_o_t(dcache_req_o_t),
     .NumPorts(NumPorts),
     .NrHwPrefetchers(NrHwPrefetchers),
     .axi_ar_chan_t(axi_ar_chan_t),
     .axi_aw_chan_t(axi_aw_chan_t),
     .axi_w_chan_t(axi_w_chan_t),
     .axi_b_chan_t(axi_b_chan_t),
     .axi_r_chan_t(axi_r_chan_t),
     .noc_req_t(noc_req_t),
     .noc_resp_t(noc_resp_t),
     .cmo_req_t(cmo_req_t),
     .cmo_rsp_t(cmo_rsp_t)
   ) i_hpdcache_subsystem (
     .clk_i(clk_i),
     .rst_ni(rst_ni),
     .noc_req_o(noc_req_o),
     .noc_resp_i(noc_resp_i),
     .icache_en_i(icache_en_i),
     .icache_flush_i(icache_flush_i),
     .icache_miss_o(icache_miss_o),
     .icache_areq_i(icache_areq_i),
     .icache_areq_o(icache_areq_o),
     .icache_dreq_i(icache_dreq_i),
     .icache_dreq_o(icache_dreq_o),
     .dcache_enable_i(dcache_enable_i),
     .dcache_flush_i(dcache_flush_i),
     .dcache_flush_ack_o(dcache_flush_ack_o),
     .dcache_miss_o(dcache_miss_o),
     .dcache_amo_req_i(dcache_amo_req_i),
     .dcache_amo_resp_o(dcache_amo_resp_o),
     .dcache_cmo_req_i(dcache_cmo_req_i),
     .dcache_cmo_resp_o(dcache_cmo_resp_o),
     .dcache_req_ports_i(dcache_req_ports_i),
     .dcache_req_ports_o(dcache_req_ports_o),
     .wbuffer_empty_o(wbuffer_empty_o),
     .wbuffer_not_ni_o(wbuffer_not_ni_o),
     .hwpf_base_set_i(hwpf_base_set_i),
     .hwpf_base_i(hwpf_base_i),
     .hwpf_base_o(hwpf_base_o),
     .hwpf_param_set_i(hwpf_param_set_i),
     .hwpf_param_i(hwpf_param_i),
     .hwpf_param_o(hwpf_param_o),
     .hwpf_throttle_set_i(hwpf_throttle_set_i),
     .hwpf_throttle_i(hwpf_throttle_i),
     .hwpf_throttle_o(hwpf_throttle_o),
     .hwpf_status_o(hwpf_status_o)
   );
endmodule
