// Copyright 2020 OpenHW Group
// Copyright 2020 Datum Technology Corporation
// Copyright 2020 Silicon Labs, Inc.
//
// Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     https://solderpad.org/licenses/
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


`ifndef __UVMA_PMA_CNTXT_SV__
`define __UVMA_PMA_CNTXT_SV__

/**
 * Object encapsulating all state variables for all PMA agent
 * (uvma_pma_agent_c) components.
 *
 * Note that the PMA Agent does not have a signal interface however the cntxt
 * is included to satisfy the base classes for uvma agents in core-v-verif
 */
class uvma_pma_cntxt_c extends uvm_object;

   `uvm_object_utils_begin(uvma_pma_cntxt_c)
   `uvm_object_utils_end

   extern function new(string name="uvma_pma_cntxt");

endclass : uvma_pma_cntxt_c


`pragma protect begin


function uvma_pma_cntxt_c::new(string name="uvma_pma_cntxt");

   super.new(name);

endfunction : new

`pragma protect end


`endif // __UVMA_PMA_CNTXT_SV__
