// COPYRIGHT HEADER


`ifndef __UVMA_RESET_MACROS_SV__
`define __UVMA_RESET_MACROS_SV__





`endif // __UVMA_RESET_MACROS_SV__
