// COPYRIGHT HEADER


`ifndef __UVMA_DEBUG_CONSTANTS_SV__
`define __UVMA_DEBUG_CONSTANTS_SV__





`endif // __UVMA_DEBUG_CONSTANTS_SV__
