/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the “License”); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File:   ariane_axi_pkg.sv
 * Author: Florian Zaruba <zarubaf@iis.ee.ethz.ch>
 * Date:   17.8.2018
 *
 * Description: Contains Ariane's AXI ports, does not contain user ports
 */

`include "axi/typedef.svh"

package ariane_axi;

    // used in axi_adapter.sv
    typedef enum logic { SINGLE_REQ, CACHE_LINE_REQ } ad_req_t;

    localparam UserWidth = 1;
    localparam AddrWidth = 64;
    localparam DataWidth = 64;
    localparam StrbWidth = DataWidth / 8;

    typedef logic [ariane_soc::IdWidth-1:0]      id_t;
    typedef logic [ariane_soc::IdWidthSlave-1:0] id_slv_t;
    typedef logic [AddrWidth-1:0] addr_t;
    typedef logic [DataWidth-1:0] data_t;
    typedef logic [StrbWidth-1:0] strb_t;
    typedef logic [UserWidth-1:0] user_t;

    `AXI_TYPEDEF_AW_CHAN_T ( aw_chan_t,     addr_t, id_t,       user_t )
    `AXI_TYPEDEF_AW_CHAN_T ( aw_chan_slv_t, addr_t, id_slv_t,   user_t )
    `AXI_TYPEDEF_W_CHAN_T  (  w_chan_t,     data_t, strb_t,     user_t )
    `AXI_TYPEDEF_B_CHAN_T  (  b_chan_t,             id_t,       user_t )
    `AXI_TYPEDEF_B_CHAN_T  (  b_chan_slv_t,         id_slv_t,   user_t )
    `AXI_TYPEDEF_AR_CHAN_T ( ar_chan_t,     addr_t, id_t,       user_t )
    `AXI_TYPEDEF_AR_CHAN_T ( ar_chan_slv_t, addr_t, id_slv_t,   user_t )
    `AXI_TYPEDEF_R_CHAN_T  (  r_chan_t,     data_t, id_t,       user_t )
    `AXI_TYPEDEF_R_CHAN_T  (  r_chan_slv_t, data_t, id_slv_t,   user_t )

    `AXI_TYPEDEF_REQ_T  ( req_t, aw_chan_t, w_chan_t, ar_chan_t )
    `AXI_TYPEDEF_RESP_T ( resp_t, b_chan_t, r_chan_t            )

    `AXI_TYPEDEF_REQ_T  ( req_slv_t, aw_chan_slv_t, w_chan_t,    ar_chan_slv_t )
    `AXI_TYPEDEF_RESP_T ( resp_slv_t, b_chan_slv_t, r_chan_slv_t               )


//    // AW Channel
//    typedef struct packed {
//        id_t              id;
//        addr_t            addr;
//        axi_pkg::len_t    len;
//        axi_pkg::size_t   size;
//        axi_pkg::burst_t  burst;
//        logic             lock;
//        axi_pkg::cache_t  cache;
//        axi_pkg::prot_t   prot;
//        axi_pkg::qos_t    qos;
//        axi_pkg::region_t region;
//        axi_pkg::atop_t   atop;
//    } aw_chan_t;
//
//    // AW Channel - Slave
//    typedef struct packed {
//        id_slv_t          id;
//        addr_t            addr;
//        axi_pkg::len_t    len;
//        axi_pkg::size_t   size;
//        axi_pkg::burst_t  burst;
//        logic             lock;
//        axi_pkg::cache_t  cache;
//        axi_pkg::prot_t   prot;
//        axi_pkg::qos_t    qos;
//        axi_pkg::region_t region;
//        axi_pkg::atop_t   atop;
//    } aw_chan_slv_t;
//
//    // W Channel - AXI4 doesn't define a wid
//    typedef struct packed {
//        data_t data;
//        strb_t strb;
//        logic  last;
//    } w_chan_t;
//
//    // B Channel
//    typedef struct packed {
//        id_t            id;
//        axi_pkg::resp_t resp;
//    } b_chan_t;
//
//    // B Channel - Slave
//    typedef struct packed {
//        id_slv_t        id;
//        axi_pkg::resp_t resp;
//    } b_chan_slv_t;
//
//    // AR Channel
//    typedef struct packed {
//        id_t             id;
//        addr_t            addr;
//        axi_pkg::len_t    len;
//        axi_pkg::size_t   size;
//        axi_pkg::burst_t  burst;
//        logic             lock;
//        axi_pkg::cache_t  cache;
//        axi_pkg::prot_t   prot;
//        axi_pkg::qos_t    qos;
//        axi_pkg::region_t region;
//    } ar_chan_t;
//
//    // AR Channel - Slave
//    typedef struct packed {
//        id_slv_t          id;
//        addr_t            addr;
//        axi_pkg::len_t    len;
//        axi_pkg::size_t   size;
//        axi_pkg::burst_t  burst;
//        logic             lock;
//        axi_pkg::cache_t  cache;
//        axi_pkg::prot_t   prot;
//        axi_pkg::qos_t    qos;
//        axi_pkg::region_t region;
//    } ar_chan_slv_t;
//
//    // R Channel
//    typedef struct packed {
//        id_t            id;
//        data_t          data;
//        axi_pkg::resp_t resp;
//        logic           last;
//    } r_chan_t;
//
//    // R Channel - Slave
//    typedef struct packed {
//        id_slv_t        id;
//        data_t          data;
//        axi_pkg::resp_t resp;
//        logic           last;
//    } r_chan_slv_t;
//
//    // Request/Response structs
//    typedef struct packed {
//        aw_chan_t aw;
//        logic     aw_valid;
//        w_chan_t  w;
//        logic     w_valid;
//        logic     b_ready;
//        ar_chan_t ar;
//        logic     ar_valid;
//        logic     r_ready;
//    } req_t;
//
//    typedef struct packed {
//        logic     aw_ready;
//        logic     ar_ready;
//        logic     w_ready;
//        logic     b_valid;
//        b_chan_t  b;
//        logic     r_valid;
//        r_chan_t  r;
//    } resp_t;
//
//    typedef struct packed {
//        aw_chan_slv_t aw;
//        logic         aw_valid;
//        w_chan_t      w;
//        logic         w_valid;
//        logic         b_ready;
//        ar_chan_slv_t ar;
//        logic         ar_valid;
//        logic         r_ready;
//    } req_slv_t;
//
//    typedef struct packed {
//        logic         aw_ready;
//        logic         ar_ready;
//        logic         w_ready;
//        logic         b_valid;
//        b_chan_slv_t  b;
//        logic         r_valid;
//        r_chan_slv_t  r;
//    } resp_slv_t;

endpackage
