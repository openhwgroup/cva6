/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 235;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00006874,
        64'h6469772D_6F692D67,
        64'h65720074_66696873,
        64'h2D676572_00737470,
        64'h75727265_746E6900,
        64'h746E6572_61702D74,
        64'h70757272_65746E69,
        64'h00646565_70732D74,
        64'h6E657272_75630076,
        64'h65646E2C_76637369,
        64'h72007974_69726F69,
        64'h72702D78_616D2C76,
        64'h63736972_0073656D,
        64'h616E2D67_65720064,
        64'h65646E65_7478652D,
        64'h73747075_72726574,
        64'h6E690073_65676E61,
        64'h7200656C_646E6168,
        64'h702C7875_6E696C00,
        64'h72656C6C_6F72746E,
        64'h6F632D74_70757272,
        64'h65746E69_00736C6C,
        64'h65632D74_70757272,
        64'h65746E69_23007469,
        64'h6C70732D_626C7400,
        64'h65707974_2D756D6D,
        64'h00617369_2C766373,
        64'h69720073_75746174,
        64'h73006765_72006570,
        64'h79745F65_63697665,
        64'h64007963_6E657571,
        64'h6572662D_6B636F6C,
        64'h63007963_6E657571,
        64'h6572662D_65736162,
        64'h656D6974_00687461,
        64'h702D7475_6F647473,
        64'h006C6564_6F6D0065,
        64'h6C626974_61706D6F,
        64'h6300736C_6C65632D,
        64'h657A6973_2300736C,
        64'h6C65632D_73736572,
        64'h64646123_09000000,
        64'h02000000_02000000,
        64'h02000000_04000000,
        64'h3A010000_04000000,
        64'h03000000_02000000,
        64'h30010000_04000000,
        64'h03000000_01000000,
        64'h25010000_04000000,
        64'h03000000_02000000,
        64'h14010000_04000000,
        64'h03000000_00C20100,
        64'h06010000_04000000,
        64'h03000000_80F0FA02,
        64'h4B000000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000010,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00303537_3631736E,
        64'h1B000000_08000000,
        64'h03000000_00000030,
        64'h30303030_30303140,
        64'h74726175_01000000,
        64'h02000000_006C6F72,
        64'h746E6F63_DE000000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000000_00000000,
        64'h67000000_10000000,
        64'h03000000_FFFF0000,
        64'h01000000_CA000000,
        64'h08000000_03000000,
        64'h00333130_2D677562,
        64'h65642C76_63736972,
        64'h1B000000_10000000,
        64'h03000000_00003040,
        64'h72656C6C_6F72746E,
        64'h6F632D67_75626564,
        64'h01000000_02000000,
        64'h02000000_BB000000,
        64'h04000000_03000000,
        64'h02000000_B5000000,
        64'h04000000_03000000,
        64'h02000000_FB000000,
        64'h04000000_03000000,
        64'h07000000_E8000000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000C_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h01000000_0B000000,
        64'h01000000_CA000000,
        64'h10000000_03000000,
        64'hA0000000_00000000,
        64'h03000000_00000030,
        64'h63696C70_2C766373,
        64'h69720030_2E302E31,
        64'h2D63696C_702C6576,
        64'h69666973_1B000000,
        64'h1E000000_03000000,
        64'h01000000_8F000000,
        64'h04000000_03000000,
        64'h00000000_00000000,
        64'h04000000_03000000,
        64'h00000000_30303030,
        64'h30306340_72656C6C,
        64'h6F72746E_6F632D74,
        64'h70757272_65746E69,
        64'h01000000_02000000,
        64'h006C6F72_746E6F63,
        64'hDE000000_08000000,
        64'h03000000_00000C00,
        64'h00000000_00000002,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h07000000_01000000,
        64'h03000000_01000000,
        64'hCA000000_10000000,
        64'h03000000_00000000,
        64'h30746E69_6C632C76,
        64'h63736972_1B000000,
        64'h0D000000_03000000,
        64'h00000030_30303030,
        64'h30324074_6E696C63,
        64'h01000000_C3000000,
        64'h00000000_03000000,
        64'h00007375_622D656C,
        64'h706D6973_00636F73,
        64'h2D657261_622D656E,
        64'h61697261_2C687465,
        64'h1B000000_1F000000,
        64'h03000000_02000000,
        64'h0F000000_04000000,
        64'h03000000_02000000,
        64'h00000000_04000000,
        64'h03000000_00636F73,
        64'h01000000_02000000,
        64'h00000008_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6F6D656D_5B000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6F6D656D,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h01000000_BB000000,
        64'h04000000_03000000,
        64'h01000000_B5000000,
        64'h04000000_03000000,
        64'h00006374_6E692D75,
        64'h70632C76_63736972,
        64'h1B000000_0F000000,
        64'h03000000_A0000000,
        64'h00000000_03000000,
        64'h01000000_8F000000,
        64'h04000000_03000000,
        64'h00000000_72656C6C,
        64'h6F72746E_6F632D74,
        64'h70757272_65746E69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732C76,
        64'h63736972_7C000000,
        64'h0B000000_03000000,
        64'h00007573_63616D69,
        64'h34367672_72000000,
        64'h0B000000_03000000,
        64'h00000076_63736972,
        64'h00656E61_69726120,
        64'h2C687465_1B000000,
        64'h12000000_03000000,
        64'h00000000_79616B6F,
        64'h6B000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5B000000_04000000,
        64'h03000000_80F0FA02,
        64'h4B000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787D01_38000000,
        64'h04000000_03000000,
        64'h00000000_0F000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313A3030_30303030,
        64'h30314074_7261752F,
        64'h636F732F_2C000000,
        64'h1A000000_03000000,
        64'h00006E65_736F6863,
        64'h01000000_00657261,
        64'h622D656E_61697261,
        64'h2C687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2D657261,
        64'h622D656E_61697261,
        64'h2C687465_1B000000,
        64'h14000000_03000000,
        64'h02000000_0F000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h54050000_47010000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h8C050000_38000000,
        64'hD3060000_EDFE0DD0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_0000BFF5,
        64'h10500073_03C58593,
        64'h00000597_F1402573,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00008402_07458593,
        64'h00000597_F1402573,
        64'h01F41413_0010041B
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
