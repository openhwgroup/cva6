// COPYRIGHT HEADER


`ifndef __UVME_CV32_MACROS_SV__
`define __UVME_CV32_MACROS_SV__





`endif // __UVME_CV32_MACROS_SV__
