// Author: Florian Zaruba, ETH Zurich, Robert Schilling, TU Graz
// Date: 27.04.2017
// Description: Abstract Sequence Item Class, similar to a UVM Sequence Item
//              Used as a common base class
//
// Copyright (C) 2017 ETH Zurich, University of Bologna
// All rights reserved.
//
// This code is under development and not yet released to the public.
// Until it is released, the code is under the copyright of ETH Zurich and
// the University of Bologna, and may contain confidential and/or unpublished
// work. Any reuse/redistribution is strictly forbidden without written
// permission from ETH Zurich.
//
// Bug fixes and contributions will eventually be released under the
// SolderPad open hardware license in the context of the PULP platform
// (http://www.pulp-platform.org), under the copyright of ETH Zurich and the
// University of Bologna.
//
class sequence_item;


endclass : sequence_item