package alu_sequence_pkg;


import fu_if_agent_pkg::*;
import uvm_pkg::*;

`include "uvm_macros.svh"
`include "fibonacci_sequence.svh"

endpackage
