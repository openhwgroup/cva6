/* File:   cache_ctrl.svh
 * Author: Florian Zaruba <zarubaf@ethz.ch>
 * Date:   14.10.2017
 *
 * Copyright (C) 2017 ETH Zurich, University of Bologna
 * All rights reserved.
 *
 * Description: Cache controller
 */
module cache_ctrl (
    input  logic clk_i,    // Clock
    input  logic rst_ni  // Asynchronous reset active low

);

endmodule
