// COPYRIGHT HEADER


`ifndef __UVML_SB_TDEFS_SV__
`define __UVML_SB_TDEFS_SV__





`endif // __UVML_SB_TDEFS_SV__
