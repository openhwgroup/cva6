`ifndef __UVMA_CORE_CNTRL_PKG_SV__
`define __UVMA_CORE_CNTRL_PKG_SV__

package uvma_core_cntrl_pkg;

   // Constants / Structs / Enums
   `include "uvma_core_cntrl_constants.sv"
   `include "uvma_core_cntrl_tdefs.sv"
   `include "uvma_core_cntrl_utils.sv"

endpackage : uvma_core_cntrl_pkg

`endif
