// COPYRIGHT HEADER


`ifndef __UVML_LOGS_MACROS_SV__
`define __UVML_LOGS_MACROS_SV__





`endif // __UVML_LOGS_MACROS_SV__
