// COPYRIGHT HEADER


`ifndef __UVML_TRN_MACROS_SV__
`define __UVML_TRN_MACROS_SV__





`endif // __UVML_TRN_MACROS_SV__
