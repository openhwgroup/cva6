// COPYRIGHT HEADER


`ifndef __UVMT_CV32_DUT_WRAP_SV__
`define __UVMT_CV32_DUT_WRAP_SV__


/**
 * Module wrapper for CV32 RTL DUT. All ports are SV interfaces.
 */
module uvmt_cv32_dut_wrap(
   uvma_debug_if  debug_if
);
   
   // TODO Instantiate Device Under Test (DUT)
   //      Ex: cv32_top  dut(
   //             .debug_data(debug_if.data),
   //             ...
   //          );
   
endmodule : uvmt_cv32_dut_wrap


`endif // __UVMT_CV32_DUT_WRAP_SV__
