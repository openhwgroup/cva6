// Enhanced memory for WT_NEW cache with proper miss handling
module wt_new_dcache_mem
  import ariane_pkg::*;
  import wt_cache_pkg::*;
  import wt_new_cache_pkg::*;
#(
  parameter config_pkg::cva6_cfg_t CVA6Cfg = config_pkg::cva6_cfg_empty,
  parameter int unsigned NUM_DUAL_SETS = wt_new_cache_pkg::NUM_DUAL_SETS,
  parameter wt_new_replacement_e REPLACEMENT_POLICY = wt_new_replacement_e'(
    REPL_ROUND_ROBIN),
  parameter wt_new_flush_policy_e FLUSH_POLICY = wt_new_flush_policy_e'(
    FLUSH_ON_SWITCH),
  parameter wt_new_b_ctrl_e B_CTRL = wt_new_b_ctrl_e'(B_CTRL_ENABLE),
  parameter type axi_req_t = logic,
  parameter type axi_rsp_t = logic
) (
  input  logic clk_i,
  input  logic rst_ni,

  // Flush dual sets when switching controllers
  input  logic flush_dual_i,

  // Controller A interface (set associative like WT cache)
  input  logic                        a_req_i,
  input  logic [CVA6Cfg.DCACHE_INDEX_WIDTH-1:0] a_index_i,
  input  logic [CVA6Cfg.DCACHE_TAG_WIDTH-1:0]   a_tag_i,
  input  logic                        a_we_i,
  input  logic [CVA6Cfg.DCACHE_LINE_WIDTH-1:0]  a_wdata_i,
  output logic [CVA6Cfg.DCACHE_LINE_WIDTH-1:0]  a_rdata_o,
  output logic                        a_hit_o,

  // Controller B interface (fully associative over dual sets)
  input  logic                        b_req_i,
  input  logic [CVA6Cfg.PLEN-1:0]     b_addr_i,
  input  logic                        b_we_i,
  input  logic [CVA6Cfg.DCACHE_LINE_WIDTH-1:0]  b_wdata_i,
  output logic [CVA6Cfg.DCACHE_LINE_WIDTH-1:0]  b_rdata_o,
  output logic                        b_hit_o,

  // Memory interface for miss handling
  output axi_req_t                    axi_data_req_o,
  input  axi_rsp_t                    axi_data_rsp_i,

  // Monitoring counters
  output logic [63:0]                 hit_count_o,
  output logic [63:0]                 miss_count_o
);

  localparam int unsigned NUM_SETS = CVA6Cfg.DCACHE_NUM_WORDS;
  localparam int unsigned ASSOC    = CVA6Cfg.DCACHE_SET_ASSOC;

  // Split memory into regular and dual-addressable sets
  localparam int unsigned NUM_REG_SETS = NUM_SETS - NUM_DUAL_SETS;

  // Cache FSM states for miss handling
  typedef enum logic [2:0] {
    IDLE,
    MISS_WAIT_GNT,
    MISS_WAIT_RESP,
    MISS_REFILL
  } cache_state_e;

  // Miss Status Holding Register (MSHR)
  typedef struct packed {
    logic                                valid;
    logic                                we;
    logic [CVA6Cfg.PLEN-1:0]            addr;
    logic [CVA6Cfg.DCACHE_LINE_WIDTH-1:0] wdata;
    logic                                is_ctrl_a;
    logic [CVA6Cfg.DCACHE_INDEX_WIDTH-1:0] index;
    logic [CVA6Cfg.DCACHE_TAG_WIDTH-1:0]   tag;
    logic [$clog2(ASSOC)-1:0]            way;
  } mshr_t;

  // Tag and data arrays
  logic [CVA6Cfg.DCACHE_TAG_WIDTH-1:0] tag_mem[NUM_SETS-1:0][ASSOC-1:0];
  logic [CVA6Cfg.DCACHE_LINE_WIDTH-1:0] data_mem[NUM_SETS-1:0][ASSOC-1:0];
  logic [ASSOC-1:0]                     valid_mem[NUM_SETS-1:0];
  logic [ASSOC-1:0]                     dirty_mem[NUM_SETS-1:0];

  // Replacement state
  logic [$clog2(NUM_DUAL_SETS)-1:0] b_repl_ptr;
  logic [CVA6Cfg.DCACHE_SET_ASSOC-1:0] a_lru_q[NUM_REG_SETS-1:0];

  // FSM state
  cache_state_e state_q, state_d;
  mshr_t mshr_q, mshr_d;

  // Memory interface signals
  logic mem_req_valid;
  logic [CVA6Cfg.PLEN-1:0] mem_req_addr;
  logic mem_req_we;
  logic [CVA6Cfg.DCACHE_LINE_WIDTH-1:0] mem_req_wdata;
  logic mem_gnt;
  logic mem_valid;
  logic [CVA6Cfg.DCACHE_LINE_WIDTH-1:0] mem_rdata;

  // Cache operation signals
  logic a_hit, b_hit_int;
  logic [CVA6Cfg.DCACHE_LINE_WIDTH-1:0] a_rdata_int, b_rdata_int;
  logic [$clog2(ASSOC)-1:0] a_hit_way, b_hit_way;
  logic [$clog2(ASSOC)-1:0] a_alloc_way;

  // Statistics counters
  logic [63:0] hit_count;
  logic [63:0] miss_count;

  // ===========================
  // Replacement Policy Logic
  // ===========================

  // Round-robin for Controller B dual sets
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      b_repl_ptr <= '0;
    end else if (b_req_i && !b_hit_int && B_CTRL == B_CTRL_ENABLE && state_q == IDLE) begin
      case (REPLACEMENT_POLICY)
        REPL_ROUND_ROBIN: b_repl_ptr <= (b_repl_ptr + 1) % NUM_DUAL_SETS;
        REPL_RANDOM: b_repl_ptr <= {$random} % NUM_DUAL_SETS;
        default: b_repl_ptr <= (b_repl_ptr + 1) % NUM_DUAL_SETS;
      endcase
    end
  end

  // LRU for Controller A regular sets
  function automatic logic [$clog2(ASSOC)-1:0] get_lru_way(
    input logic [ASSOC-1:0] valid,
    input logic [ASSOC-1:0] lru_state
  );
    // Find first invalid way, or LRU way if all valid
    for (int i = 0; i < ASSOC; i++) begin
      if (!valid[i]) return i;
    end
    // All ways valid, return LRU (simplified - just round robin)
    for (int i = 0; i < ASSOC; i++) begin
      if (lru_state[i]) return i;
    end
    return 0;
  endfunction

  // Update LRU on access
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      a_lru_q <= '{default: '0};
    end else if (a_req_i && a_hit && a_index_i < NUM_REG_SETS) begin
      // Update LRU - move accessed way to MRU position (only for regular sets)
      a_lru_q[a_index_i] <= (a_lru_q[a_index_i] + 1) % ASSOC;
    end
  end

  // ===========================
  // Cache Tag/Data Access Logic
  // ===========================

  // Controller A tag comparison (all ways)
  always_comb begin
    a_hit = 1'b0;
    a_hit_way = '0;
    a_rdata_int = '0;
    if (a_index_i < NUM_REG_SETS) begin
      a_alloc_way = get_lru_way(valid_mem[a_index_i], a_lru_q[a_index_i]);
    end else begin
      a_alloc_way = 0; // For dual sets, Controller A only uses way 0
    end
    
    for (int way = 0; way < ASSOC; way++) begin
      if (valid_mem[a_index_i][way] && 
          tag_mem[a_index_i][way] == a_tag_i) begin
        a_hit = 1'b1;
        a_hit_way = way;
        a_rdata_int = data_mem[a_index_i][way];
        break;
      end
    end
  end

  // Controller B tag comparison (dual sets only)
  always_comb begin
    b_hit_int = 1'b0;
    b_hit_way = '0;
    b_rdata_int = '0;
    
    if (B_CTRL == B_CTRL_ENABLE) begin
      // Hash-based lookup optimization for PSEUDO_LRU
      if (REPLACEMENT_POLICY == REPL_PSEUDO_LRU) begin
        int lookup_idx = NUM_REG_SETS + (b_addr_i[3:2] % NUM_DUAL_SETS);
        if (valid_mem[lookup_idx][0] &&
            tag_mem[lookup_idx][0] == b_addr_i[CVA6Cfg.DCACHE_TAG_WIDTH+CVA6Cfg.DCACHE_INDEX_WIDTH-1:CVA6Cfg.DCACHE_INDEX_WIDTH]) begin
          b_hit_int = 1'b1;
          b_hit_way = 0;
          b_rdata_int = data_mem[lookup_idx][0];
        end
      end
      
      // Linear search if hash miss or other policies
      if (!b_hit_int) begin
        for (int s = 0; s < NUM_DUAL_SETS; s++) begin
          int idx = NUM_REG_SETS + s;
          if (valid_mem[idx][0] &&
              tag_mem[idx][0] == b_addr_i[CVA6Cfg.DCACHE_TAG_WIDTH+CVA6Cfg.DCACHE_INDEX_WIDTH-1:CVA6Cfg.DCACHE_INDEX_WIDTH]) begin
            b_hit_int = 1'b1;
            b_hit_way = 0;
            b_rdata_int = data_mem[idx][0];
            break;
          end
        end
      end
    end
  end

  // ===========================
  // Miss Handling FSM
  // ===========================

  always_comb begin
    state_d = state_q;
    mshr_d = mshr_q;
    
    mem_req_valid = 1'b0;
    mem_req_addr = '0;
    mem_req_we = 1'b0;
    mem_req_wdata = '0;

    case (state_q)
      IDLE: begin
        // Check for cache misses
        if (a_req_i && !a_hit && !a_we_i) begin
          // Controller A read miss
          state_d = MISS_WAIT_GNT;
          mshr_d.valid = 1'b1;
          mshr_d.we = a_we_i;
          mshr_d.addr = {a_tag_i, a_index_i, {CVA6Cfg.DCACHE_OFFSET_WIDTH{1'b0}}};
          mshr_d.wdata = a_wdata_i;
          mshr_d.is_ctrl_a = 1'b1;
          mshr_d.index = a_index_i;
          mshr_d.tag = a_tag_i;
          if (a_index_i < NUM_REG_SETS) begin
            mshr_d.way = get_lru_way(valid_mem[a_index_i], a_lru_q[a_index_i]);
          end else begin
            mshr_d.way = 0; // For dual sets, Controller A only uses way 0
          end
        end else if (b_req_i && !b_hit_int && !b_we_i && B_CTRL == B_CTRL_ENABLE) begin
          // Controller B read miss
          state_d = MISS_WAIT_GNT;
          mshr_d.valid = 1'b1;
          mshr_d.we = b_we_i;
          mshr_d.addr = {b_addr_i[CVA6Cfg.PLEN-1:CVA6Cfg.DCACHE_OFFSET_WIDTH], {CVA6Cfg.DCACHE_OFFSET_WIDTH{1'b0}}};
          mshr_d.wdata = b_wdata_i;
          mshr_d.is_ctrl_a = 1'b0;
          mshr_d.index = NUM_REG_SETS + b_repl_ptr;
          mshr_d.tag = b_addr_i[CVA6Cfg.DCACHE_TAG_WIDTH+CVA6Cfg.DCACHE_INDEX_WIDTH-1:CVA6Cfg.DCACHE_INDEX_WIDTH];
          mshr_d.way = 0; // Controller B uses way 0 only
        end
      end

      MISS_WAIT_GNT: begin
        mem_req_valid = 1'b1;
        mem_req_addr = mshr_q.addr;
        mem_req_we = 1'b0; // Read from memory
        
        if (mem_gnt) begin
          state_d = MISS_WAIT_RESP;
        end
      end

      MISS_WAIT_RESP: begin
        if (mem_valid) begin
          state_d = MISS_REFILL;
        end
      end

      MISS_REFILL: begin
        // Cache line refill completed in next cycle
        state_d = IDLE;
        mshr_d.valid = 1'b0;
      end

      default: state_d = IDLE;
    endcase
  end

  // ===========================
  // Cache Array Updates
  // ===========================

  // Flush dual sets on controller switch
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      valid_mem <= '{default: '0};
      dirty_mem <= '{default: '0};
    end else if (flush_dual_i && FLUSH_POLICY == FLUSH_ON_SWITCH) begin
      // Flush only dual sets
      valid_mem[NUM_REG_SETS+:NUM_DUAL_SETS] <= '{default: '0};
      dirty_mem[NUM_REG_SETS+:NUM_DUAL_SETS] <= '{default: '0};
    end else begin
      // Normal cache operations
      
      // Controller A write operations
      if (a_req_i && a_we_i && state_q == IDLE) begin
        if (a_hit) begin
          // Write hit - update existing line
          data_mem[a_index_i][a_hit_way] <= a_wdata_i;
          dirty_mem[a_index_i][a_hit_way] <= 1'b1;
        end else begin
          // Write miss - allocate new line (write-allocate)
          tag_mem[a_index_i][a_alloc_way] <= a_tag_i;
          data_mem[a_index_i][a_alloc_way] <= a_wdata_i;
          valid_mem[a_index_i][a_alloc_way] <= 1'b1;
          dirty_mem[a_index_i][a_alloc_way] <= 1'b1;
        end
      end

      // Controller B write operations
      if (b_req_i && b_we_i && B_CTRL == B_CTRL_ENABLE && state_q == IDLE) begin
        if (b_hit_int) begin
          // Write hit - find the hitting way
          for (int s = 0; s < NUM_DUAL_SETS; s++) begin
            int idx = NUM_REG_SETS + s;
            if (valid_mem[idx][0] &&
                tag_mem[idx][0] == b_addr_i[CVA6Cfg.DCACHE_TAG_WIDTH+CVA6Cfg.DCACHE_INDEX_WIDTH-1:CVA6Cfg.DCACHE_INDEX_WIDTH]) begin
              data_mem[idx][0] = b_wdata_i;
              dirty_mem[idx][0] = 1'b1;
              break;
            end
          end
        end else begin
          // Write miss - allocate using replacement policy
          int alloc_idx = NUM_REG_SETS + b_repl_ptr;
          tag_mem[alloc_idx][0] <= b_addr_i[CVA6Cfg.DCACHE_TAG_WIDTH+CVA6Cfg.DCACHE_INDEX_WIDTH-1:CVA6Cfg.DCACHE_INDEX_WIDTH];
          data_mem[alloc_idx][0] <= b_wdata_i;
          valid_mem[alloc_idx][0] <= 1'b1;
          dirty_mem[alloc_idx][0] <= 1'b1;
        end
      end

      // Cache line refill from memory
      if (state_q == MISS_REFILL && mem_valid) begin
        if (mshr_q.is_ctrl_a) begin
          tag_mem[mshr_q.index][mshr_q.way] <= mshr_q.tag;
          data_mem[mshr_q.index][mshr_q.way] <= mem_rdata;
          valid_mem[mshr_q.index][mshr_q.way] <= 1'b1;
          dirty_mem[mshr_q.index][mshr_q.way] <= 1'b0;
        end else begin
          tag_mem[mshr_q.index][mshr_q.way] <= mshr_q.tag;
          data_mem[mshr_q.index][mshr_q.way] <= mem_rdata;
          valid_mem[mshr_q.index][mshr_q.way] <= 1'b1;
          dirty_mem[mshr_q.index][mshr_q.way] <= 1'b0;
        end
      end
    end
  end

  // ===========================
  // Output Assignment
  // ===========================

  always_comb begin
    // Controller A outputs
    if (state_q == MISS_REFILL && mshr_q.is_ctrl_a && mem_valid) begin
      a_rdata_o = mem_rdata;
      a_hit_o = 1'b1;
    end else if (state_q != IDLE && mshr_q.is_ctrl_a) begin
      // During miss handling, report miss
      a_rdata_o = '0;
      a_hit_o = 1'b0;
    end else begin
      a_rdata_o = a_hit ? a_rdata_int : '0;
      a_hit_o = a_hit && (state_q == IDLE);
    end

    // Controller B outputs  
    if (state_q == MISS_REFILL && !mshr_q.is_ctrl_a && mem_valid) begin
      b_rdata_o = mem_rdata;
      b_hit_o = 1'b1;
    end else if (state_q != IDLE && !mshr_q.is_ctrl_a) begin
      // During miss handling, report miss
      b_rdata_o = '0;
      b_hit_o = 1'b0;
    end else if (b_we_i) begin
      // Write operations always "hit" (write-allocate)
      b_rdata_o = '0;
      b_hit_o = 1'b1;
    end else begin
      b_rdata_o = b_hit_int ? b_rdata_int : '0;
      b_hit_o = b_hit_int && (state_q == IDLE);
    end
  end

  // Count hits and misses
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      hit_count <= '0;
      miss_count <= '0;
    end else begin
      if (a_req_i && !a_we_i) begin
        if (a_hit || (state_q == MISS_REFILL && mshr_q.is_ctrl_a)) hit_count <= hit_count + 1;
        else if (state_q == IDLE) miss_count <= miss_count + 1;
      end
      if (b_req_i && !b_we_i && B_CTRL == B_CTRL_ENABLE) begin
        if (b_hit_int || (state_q == MISS_REFILL && !mshr_q.is_ctrl_a)) hit_count <= hit_count + 1;
        else if (state_q == IDLE) miss_count <= miss_count + 1;
      end
    end
  end

  // FSM state register
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      state_q <= IDLE;
      mshr_q <= '0;
    end else begin
      state_q <= state_d;
      mshr_q <= mshr_d;
    end
  end

  assign hit_count_o = hit_count;
  assign miss_count_o = miss_count;

  // ===========================
  // AXI Interface for Memory
  // ===========================

  // Simplified AXI interface - would need proper AXI adapter in real implementation
  assign axi_data_req_o.aw_valid = mem_req_valid && mem_req_we;
  assign axi_data_req_o.aw.addr = mem_req_addr;
  assign axi_data_req_o.aw.id = '0;
  assign axi_data_req_o.aw.len = '0;
  assign axi_data_req_o.aw.size = 3'b011; // 8 bytes
  assign axi_data_req_o.aw.burst = 2'b01; // INCR
  assign axi_data_req_o.aw.lock = '0;
  assign axi_data_req_o.aw.cache = '0;
  assign axi_data_req_o.aw.prot = '0;
  assign axi_data_req_o.aw.qos = '0;
  assign axi_data_req_o.aw.region = '0;
  assign axi_data_req_o.aw.atop = '0;
  assign axi_data_req_o.aw.user = '0;

  assign axi_data_req_o.w_valid = mem_req_valid && mem_req_we;
  assign axi_data_req_o.w.data = mem_req_wdata;
  assign axi_data_req_o.w.strb = '1;
  assign axi_data_req_o.w.last = 1'b1;
  assign axi_data_req_o.w.user = '0;

  assign axi_data_req_o.ar_valid = mem_req_valid && !mem_req_we;
  assign axi_data_req_o.ar.addr = mem_req_addr;
  assign axi_data_req_o.ar.id = '0;
  assign axi_data_req_o.ar.len = '0;
  assign axi_data_req_o.ar.size = 3'b011; // 8 bytes
  assign axi_data_req_o.ar.burst = 2'b01; // INCR
  assign axi_data_req_o.ar.lock = '0;
  assign axi_data_req_o.ar.cache = '0;
  assign axi_data_req_o.ar.prot = '0;
  assign axi_data_req_o.ar.qos = '0;
  assign axi_data_req_o.ar.region = '0;
  assign axi_data_req_o.ar.user = '0;

  assign axi_data_req_o.r_ready = 1'b1;
  assign axi_data_req_o.b_ready = 1'b1;

  assign mem_gnt = mem_req_we ? (axi_data_rsp_i.aw_ready && axi_data_rsp_i.w_ready) : 
                                axi_data_rsp_i.ar_ready;
  assign mem_valid = mem_req_we ? axi_data_rsp_i.b_valid : axi_data_rsp_i.r_valid;
  assign mem_rdata = axi_data_rsp_i.r.data;
endmodule
