/*
 *
 * Copyright (c) 2005-2020 Imperas Software Ltd., All Rights Reserved.
 *
 * THIS SOFTWARE CONTAINS CONFIDENTIAL INFORMATION AND TRADE SECRETS
 * OF IMPERAS SOFTWARE LTD. USE, DISCLOSURE, OR REPRODUCTION IS PROHIBITED
 * EXCEPT AS MAY BE PROVIDED FOR IN A WRITTEN AGREEMENT WITH
 * IMPERAS SOFTWARE LTD.
 *
 */

`ifndef __INCL_TYPEDEFS_SV
`define __INCL_TYPEDEFS_SV

//
// Address label monitor type
//
typedef struct {
    int addr;
    int enable;
} watchT;

typedef int unsigned Uns32;

`endif