// COPYRIGHT HEADER


`ifndef __UVMT_CV32_CONSTANTS_SV__
`define __UVMT_CV32_CONSTANTS_SV__





`endif // __UVMT_CV32_CONSTANTS_SV__
