// Copyright 2020 OpenHW Group
// Copyright 2020 Datum Technology Corporation
// Copyright 2020 Silicon Labs, Inc.
//
// Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     https://solderpad.org/licenses/
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


`ifndef __UVMA_FENCEI_TDEFS_SV__
`define __UVMA_FENCEI_TDEFS_SV__

typedef enum {
   UVMA_FENCEI_DRV_ACK_MODE_CONSTANT,
   UVMA_FENCEI_DRV_ACK_MODE_FIXED_LATENCY,
   UVMA_FENCEI_DRV_ACK_MODE_RANDOM_LATENCY
} uvma_fencei_drv_ack_enum;

typedef enum {
   UVMA_FENCEI_RESET_STATE_PRE_RESET ,
   UVMA_FENCEI_RESET_STATE_IN_RESET  ,
   UVMA_FENCEI_RESET_STATE_POST_RESET
} uvma_fencei_reset_state_enum;


`endif // __UVMA_FENCEI_TDEFS_SV__
