// 
// Copyright 2020 OpenHW Group
// Copyright 2020 Datum Technology Corporation
// 
// Licensed under the Solderpad Hardware License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// 
//     https://solderpad.org/licenses/
// 
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// 


`ifndef __UVML_HRTBT_CONSTANTS_SV__
`define __UVML_HRTBT_CONSTANTS_SV__


<<<<<<< HEAD
const int unsigned  uvml_hrtbt_default_startup_timeout  = 10_000;
const int unsigned  uvml_hrtbt_default_heartbeat_period = 20_000;
const int unsigned  uvml_hrtbt_default_refresh_period   =  5_000;
=======
const int unsigned  uvm_hrtbt_default_startup_timeout  = 10_000;
const int unsigned  uvm_hrtbt_default_heartbeat_period = 20_000;
const int unsigned  uvm_hrtbt_default_refresh_period   =  5_000;
>>>>>>> 3f88a4d93395bc9a977a691a2503368f7eda98dc


`endif // __UVML_HRTBT_CONSTANTS_SV__
