/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the “License”); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 211;

    const logic [RomSize-1:0][63:0] mem = {
        64'h006b,
        64'h636f6c63_00737470,
        64'h75727265_746e6900,
        64'h746e6572_61702d74,
        64'h70757272_65746e69,
        64'h00766564_6e2c7663,
        64'h73697200_79746972,
        64'h6f697270_2d78616d,
        64'h2c766373_69720073,
        64'h656d616e_2d676572,
        64'h00646564_6e657478,
        64'h652d7374_70757272,
        64'h65746e69_00736567,
        64'h6e617200_656c646e,
        64'h6168702c_78756e69,
        64'h6c007265_6c6c6f72,
        64'h746e6f63_2d747075,
        64'h72726574_6e690073,
        64'h6c6c6563_2d747075,
        64'h72726574_6e692300,
        64'h79636e65_75716572,
        64'h662d6b63_6f6c6300,
        64'h65707974_2d756d6d,
        64'h00617369_2c766373,
        64'h69720073_75746174,
        64'h73006765_72006570,
        64'h79745f65_63697665,
        64'h64007963_6e657571,
        64'h6572662d_65736162,
        64'h656d6974_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h80f0fa02_0c010000,
        64'h04000000_03000000,
        64'h02000000_01000000,
        64'h00000000_01010000,
        64'h0c000000_03000000,
        64'h02000000_f0000000,
        64'h04000000_03000000,
        64'h00000100_00000000,
        64'h00000010_00000000,
        64'h4b000000_10000000,
        64'h03000000_00000000,
        64'h612e3230_2e312d65,
        64'h74696c74_7261752d,
        64'h6978612c_786e6c78,
        64'h1b000000_19000000,
        64'h03000000_00000030,
        64'h30303030_30303140,
        64'h74726175_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_c8000000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000000_00000000,
        64'h4b000000_10000000,
        64'h03000000_ffff0000,
        64'h01000000_b4000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00003040,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h02000000_a5000000,
        64'h04000000_03000000,
        64'h02000000_9f000000,
        64'h04000000_03000000,
        64'h35000000_e5000000,
        64'h04000000_03000000,
        64'h07000000_d2000000,
        64'h04000000_03000000,
        64'h006c6f72_746e6f63,
        64'hc8000000_08000000,
        64'h03000000_00000004,
        64'h00000000_0000000c,
        64'h00000000_4b000000,
        64'h10000000_03000000,
        64'h09000000_01000000,
        64'h0b000000_01000000,
        64'hb4000000_10000000,
        64'h03000000_8a000000,
        64'h00000000_03000000,
        64'h00306369_6c702c76,
        64'h63736972_1b000000,
        64'h0c000000_03000000,
        64'h01000000_79000000,
        64'h04000000_03000000,
        64'h00000000_30303030,
        64'h30306340_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_02000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h4b000000_10000000,
        64'h03000000_07000000,
        64'h01000000_03000000,
        64'h01000000_b4000000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'had000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_00000002,
        64'h00000000_00000080,
        64'h00000000_4b000000,
        64'h10000000_03000000,
        64'h00007972_6f6d656d,
        64'h3f000000_07000000,
        64'h03000000_00303030,
        64'h30303030_38407972,
        64'h6f6d656d_01000000,
        64'h02000000_02000000,
        64'h02000000_01000000,
        64'ha5000000_04000000,
        64'h03000000_01000000,
        64'h9f000000_04000000,
        64'h03000000_00006374,
        64'h6e692d75_70632c76,
        64'h63736972_1b000000,
        64'h0f000000_03000000,
        64'h8a000000_00000000,
        64'h03000000_01000000,
        64'h79000000_04000000,
        64'h03000000_00000000,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h80f0fa02_69000000,
        64'h04000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_60000000,
        64'h0b000000_03000000,
        64'h00636d69_34367672,
        64'h56000000_08000000,
        64'h03000000_00000076,
        64'h63736972_1b000000,
        64'h06000000_03000000,
        64'h00000000_79616b6f,
        64'h4f000000_05000000,
        64'h03000000_00000000,
        64'h4b000000_04000000,
        64'h03000000_00757063,
        64'h3f000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_2c000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hc8040000_12010000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h00050000_38000000,
        64'h12060000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_0000bff5,
        64'h10500073_03c58593,
        64'h00000597_f1402573,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00008402_07458593,
        64'h00000597_f1402573,
        64'h01f41413_0010041b
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    assign rdata_o = mem[addr_q];
endmodule
