module axi_crossbar_wrap (
AXI_BUS.Slave slave0_if, slave1_if, slave2_if, slave3_if,
AXI_BUS.Master master0_if, master1_if, master2_if,
input clk_i, rst_ni
);
  
axi_crossbar_0 your_instance_name (
  .aclk(clk_i),                   // input wire aclk
  .aresetn(rst_ni),             // input wire aresetn
  .s_axi_awid({slave3_if.aw_id,slave2_if.aw_id,slave1_if.aw_id,slave0_if.aw_id}),
  .s_axi_awaddr({slave3_if.aw_addr,slave2_if.aw_addr,slave1_if.aw_addr,slave0_if.aw_addr}),
  .s_axi_awlen({slave3_if.aw_len,slave2_if.aw_len,slave1_if.aw_len,slave0_if.aw_len}),
  .s_axi_awsize({slave3_if.aw_size,slave2_if.aw_size,slave1_if.aw_size,slave0_if.aw_size}),
  .s_axi_awburst({slave3_if.aw_burst,slave2_if.aw_burst,slave1_if.aw_burst,slave0_if.aw_burst}),
  .s_axi_awlock({slave3_if.aw_lock,slave2_if.aw_lock,slave1_if.aw_lock,slave0_if.aw_lock}),
  .s_axi_awcache({slave3_if.aw_cache,slave2_if.aw_cache,slave1_if.aw_cache,slave0_if.aw_cache}),
  .s_axi_awprot({slave3_if.aw_prot,slave2_if.aw_prot,slave1_if.aw_prot,slave0_if.aw_prot}),
//.s_axi_awregion({slave3_if.aw_region,slave2_if.aw_region,slave1_if.aw_region,slave0_if.aw_region}),
  .s_axi_awqos({slave3_if.aw_qos,slave2_if.aw_qos,slave1_if.aw_qos,slave0_if.aw_qos}),
  .s_axi_awuser({slave3_if.aw_user,slave2_if.aw_user,slave1_if.aw_user,slave0_if.aw_user}),
  .s_axi_awvalid({slave3_if.aw_valid,slave2_if.aw_valid,slave1_if.aw_valid,slave0_if.aw_valid}),
  .s_axi_awready({slave3_if.aw_ready,slave2_if.aw_ready,slave1_if.aw_ready,slave0_if.aw_ready}),
  .s_axi_wdata({slave3_if.w_data,slave2_if.w_data,slave1_if.w_data,slave0_if.w_data}),
  .s_axi_wstrb({slave3_if.w_strb,slave2_if.w_strb,slave1_if.w_strb,slave0_if.w_strb}),
  .s_axi_wlast({slave3_if.w_last,slave2_if.w_last,slave1_if.w_last,slave0_if.w_last}),
  .s_axi_wuser({slave3_if.w_user,slave2_if.w_user,slave1_if.w_user,slave0_if.w_user}),
  .s_axi_wvalid({slave3_if.w_valid,slave2_if.w_valid,slave1_if.w_valid,slave0_if.w_valid}),
  .s_axi_wready({slave3_if.w_ready,slave2_if.w_ready,slave1_if.w_ready,slave0_if.w_ready}),
  .s_axi_bid({slave3_if.b_id,slave2_if.b_id,slave1_if.b_id,slave0_if.b_id}),
  .s_axi_bresp({slave3_if.b_resp,slave2_if.b_resp,slave1_if.b_resp,slave0_if.b_resp}),
  .s_axi_buser({slave3_if.b_user,slave2_if.b_user,slave1_if.b_user,slave0_if.b_user}),
  .s_axi_bvalid({slave3_if.b_valid,slave2_if.b_valid,slave1_if.b_valid,slave0_if.b_valid}),
  .s_axi_bready({slave3_if.b_ready,slave2_if.b_ready,slave1_if.b_ready,slave0_if.b_ready}),
  .s_axi_arid({slave3_if.ar_id,slave2_if.ar_id,slave1_if.ar_id,slave0_if.ar_id}),
  .s_axi_araddr({slave3_if.ar_addr,slave2_if.ar_addr,slave1_if.ar_addr,slave0_if.ar_addr}),
  .s_axi_arlen({slave3_if.ar_len,slave2_if.ar_len,slave1_if.ar_len,slave0_if.ar_len}),
  .s_axi_arsize({slave3_if.ar_size,slave2_if.ar_size,slave1_if.ar_size,slave0_if.ar_size}),
  .s_axi_arburst({slave3_if.ar_burst,slave2_if.ar_burst,slave1_if.ar_burst,slave0_if.ar_burst}),
  .s_axi_arlock({slave3_if.ar_lock,slave2_if.ar_lock,slave1_if.ar_lock,slave0_if.ar_lock}),
  .s_axi_arcache({slave3_if.ar_cache,slave2_if.ar_cache,slave1_if.ar_cache,slave0_if.ar_cache}),
  .s_axi_arprot({slave3_if.ar_prot,slave2_if.ar_prot,slave1_if.ar_prot,slave0_if.ar_prot}),
//  .s_axi_arregion({slave3_if.ar_region,slave2_if.ar_region,slave1_if.ar_region,slave0_if.ar_region}),
  .s_axi_arqos({slave3_if.ar_qos,slave2_if.ar_qos,slave1_if.ar_qos,slave0_if.ar_qos}),
  .s_axi_aruser({slave3_if.ar_user,slave2_if.ar_user,slave1_if.ar_user,slave0_if.ar_user}),
  .s_axi_arvalid({slave3_if.ar_valid,slave2_if.ar_valid,slave1_if.ar_valid,slave0_if.ar_valid}),
  .s_axi_arready({slave3_if.ar_ready,slave2_if.ar_ready,slave1_if.ar_ready,slave0_if.ar_ready}),
  .s_axi_rid({slave3_if.r_id,slave2_if.r_id,slave1_if.r_id,slave0_if.r_id}),
  .s_axi_rdata({slave3_if.r_data,slave2_if.r_data,slave1_if.r_data,slave0_if.r_data}),
  .s_axi_rresp({slave3_if.r_resp,slave2_if.r_resp,slave1_if.r_resp,slave0_if.r_resp}),
  .s_axi_rlast({slave3_if.r_last,slave2_if.r_last,slave1_if.r_last,slave0_if.r_last}),
  .s_axi_ruser({slave3_if.r_user,slave2_if.r_user,slave1_if.r_user,slave0_if.r_user}),
  .s_axi_rvalid({slave3_if.r_valid,slave2_if.r_valid,slave1_if.r_valid,slave0_if.r_valid}),
  .s_axi_rready({slave3_if.r_ready,slave2_if.r_ready,slave1_if.r_ready,slave0_if.r_ready}),
    .m_axi_awvalid  ( {master2_if.aw_valid , master1_if.aw_valid , master0_if.aw_valid } ),
    .m_axi_awaddr   ( {master2_if.aw_addr  , master1_if.aw_addr  , master0_if.aw_addr  } ),
    .m_axi_awprot   ( {master2_if.aw_prot  , master1_if.aw_prot  , master0_if.aw_prot  } ),
    .m_axi_awregion ( {master2_if.aw_region, master1_if.aw_region, master0_if.aw_region} ),
    .m_axi_awlen    ( {master2_if.aw_len   , master1_if.aw_len   , master0_if.aw_len   } ),
    .m_axi_awsize   ( {master2_if.aw_size  , master1_if.aw_size  , master0_if.aw_size  } ),
    .m_axi_awburst  ( {master2_if.aw_burst , master1_if.aw_burst , master0_if.aw_burst } ),
    .m_axi_awlock   ( {master2_if.aw_lock  , master1_if.aw_lock  , master0_if.aw_lock  } ),
    .m_axi_awcache  ( {master2_if.aw_cache , master1_if.aw_cache , master0_if.aw_cache } ),
    .m_axi_awqos    ( {master2_if.aw_qos   , master1_if.aw_qos   , master0_if.aw_qos   } ),
    .m_axi_awid     ( {master2_if.aw_id    , master1_if.aw_id    , master0_if.aw_id    } ),
    .m_axi_awuser   ( {master2_if.aw_user  , master1_if.aw_user  , master0_if.aw_user  } ),
    .m_axi_awready  ( {master2_if.aw_ready , master1_if.aw_ready , master0_if.aw_ready } ),

    .m_axi_arvalid  ( {master2_if.ar_valid , master1_if.ar_valid , master0_if.ar_valid } ),
    .m_axi_araddr   ( {master2_if.ar_addr  , master1_if.ar_addr  , master0_if.ar_addr  } ),
    .m_axi_arprot   ( {master2_if.ar_prot  , master1_if.ar_prot  , master0_if.ar_prot  } ),
    .m_axi_arregion ( {master2_if.ar_region, master1_if.ar_region, master0_if.ar_region} ),
    .m_axi_arlen    ( {master2_if.ar_len   , master1_if.ar_len   , master0_if.ar_len   } ),
    .m_axi_arsize   ( {master2_if.ar_size  , master1_if.ar_size  , master0_if.ar_size  } ),
    .m_axi_arburst  ( {master2_if.ar_burst , master1_if.ar_burst , master0_if.ar_burst } ),
    .m_axi_arlock   ( {master2_if.ar_lock  , master1_if.ar_lock  , master0_if.ar_lock  } ),
    .m_axi_arcache  ( {master2_if.ar_cache , master1_if.ar_cache , master0_if.ar_cache } ),
    .m_axi_arqos    ( {master2_if.ar_qos   , master1_if.ar_qos   , master0_if.ar_qos   } ),
    .m_axi_arid     ( {master2_if.ar_id    , master1_if.ar_id    , master0_if.ar_id    } ),
    .m_axi_aruser   ( {master2_if.ar_user  , master1_if.ar_user  , master0_if.ar_user  } ),
    .m_axi_arready  ( {master2_if.ar_ready , master1_if.ar_ready , master0_if.ar_ready } ),

    .m_axi_wvalid   ( {master2_if.w_valid  , master1_if.w_valid  , master0_if.w_valid  } ),
//    .m_axi_wid      ( {master2_if.w_id     , master1_if.w_id     , master0_if.w_id     } ),
    .m_axi_wdata    ( {master2_if.w_data   , master1_if.w_data   , master0_if.w_data   } ),
    .m_axi_wstrb    ( {master2_if.w_strb   , master1_if.w_strb   , master0_if.w_strb   } ),
    .m_axi_wuser    ( {master2_if.w_user   , master1_if.w_user   , master0_if.w_user   } ),
    .m_axi_wlast    ( {master2_if.w_last   , master1_if.w_last   , master0_if.w_last   } ),
    .m_axi_wready   ( {master2_if.w_ready  , master1_if.w_ready  , master0_if.w_ready  } ),

    .m_axi_rvalid   ( {master2_if.r_valid  , master1_if.r_valid  , master0_if.r_valid  } ),
    .m_axi_rdata    ( {master2_if.r_data   , master1_if.r_data   , master0_if.r_data   } ),
    .m_axi_rresp    ( {master2_if.r_resp   , master1_if.r_resp   , master0_if.r_resp   } ),
    .m_axi_rlast    ( {master2_if.r_last   , master1_if.r_last   , master0_if.r_last   } ),
    .m_axi_rid      ( {master2_if.r_id     , master1_if.r_id     , master0_if.r_id     } ),
    .m_axi_ruser    ( {master2_if.r_user   , master1_if.r_user   , master0_if.r_user   } ),
    .m_axi_rready   ( {master2_if.r_ready  , master1_if.r_ready  , master0_if.r_ready  } ),

    .m_axi_bvalid   ( {master2_if.b_valid  , master1_if.b_valid  , master0_if.b_valid  } ),
    .m_axi_bresp    ( {master2_if.b_resp   , master1_if.b_resp   , master0_if.b_resp   } ),
    .m_axi_bid      ( {master2_if.b_id     , master1_if.b_id     , master0_if.b_id     } ),
    .m_axi_buser    ( {master2_if.b_user   , master1_if.b_user   , master0_if.b_user   } ),
    .m_axi_bready   ( {master2_if.b_ready  , master1_if.b_ready  , master0_if.b_ready  } )
);

endmodule // nasti_converter
