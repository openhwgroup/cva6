/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 236;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00006874,
        64'h61702D74_756F6474,
        64'h73006874_6469772D,
        64'h6F692D67_65720074,
        64'h66696873_2D676572,
        64'h00737470_75727265,
        64'h746E6900_746E6572,
        64'h61702D74_70757272,
        64'h65746E69_00646565,
        64'h70732D74_6E657272,
        64'h75630076_65646E2C,
        64'h76637369_72007974,
        64'h69726F69_72702D78,
        64'h616D2C76_63736972,
        64'h0073656D_616E2D67,
        64'h65720064_65646E65,
        64'h7478652D_73747075,
        64'h72726574_6E690073,
        64'h65676E61_7200656C,
        64'h646E6168_702C7875,
        64'h6E696C00_72656C6C,
        64'h6F72746E_6F632D74,
        64'h70757272_65746E69,
        64'h00736C6C_65632D74,
        64'h70757272_65746E69,
        64'h23007469_6C70732D,
        64'h626C7400_65707974,
        64'h2D756D6D_00617369,
        64'h2C766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745F65,
        64'h63697665_64007963,
        64'h6E657571_6572662D,
        64'h6B636F6C_63007963,
        64'h6E657571_6572662D,
        64'h65736162_656D6974,
        64'h006C6564_6F6D0065,
        64'h6C626974_61706D6F,
        64'h6300736C_6C65632D,
        64'h657A6973_2300736C,
        64'h6C65632D_73736572,
        64'h64646123_09000000,
        64'h02000000_02000000,
        64'h00003030_30303030,
        64'h30314074_7261752F,
        64'h636F732F_3B010000,
        64'h13000000_03000000,
        64'h00006E65_736F6863,
        64'h01000000_02000000,
        64'h02000000_04000000,
        64'h2E010000_04000000,
        64'h03000000_02000000,
        64'h24010000_04000000,
        64'h03000000_01000000,
        64'h19010000_04000000,
        64'h03000000_02000000,
        64'h08010000_04000000,
        64'h03000000_00C20100,
        64'hFA000000_04000000,
        64'h03000000_80F0FA02,
        64'h3F000000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000010,
        64'h00000000_5B000000,
        64'h10000000_03000000,
        64'h00303537_3631736E,
        64'h1B000000_08000000,
        64'h03000000_00000030,
        64'h30303030_30303140,
        64'h74726175_01000000,
        64'h02000000_006C6F72,
        64'h746E6F63_D2000000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000000_00000000,
        64'h5B000000_10000000,
        64'h03000000_FFFF0000,
        64'h01000000_BE000000,
        64'h08000000_03000000,
        64'h00333130_2D677562,
        64'h65642C76_63736972,
        64'h1B000000_10000000,
        64'h03000000_00003040,
        64'h72656C6C_6F72746E,
        64'h6F632D67_75626564,
        64'h01000000_02000000,
        64'h02000000_AF000000,
        64'h04000000_03000000,
        64'h02000000_A9000000,
        64'h04000000_03000000,
        64'h02000000_EF000000,
        64'h04000000_03000000,
        64'h07000000_DC000000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000C_00000000,
        64'h5B000000_10000000,
        64'h03000000_09000000,
        64'h01000000_0B000000,
        64'h01000000_BE000000,
        64'h10000000_03000000,
        64'h94000000_00000000,
        64'h03000000_00000030,
        64'h63696C70_2C766373,
        64'h69720030_2E302E31,
        64'h2D63696C_702C6576,
        64'h69666973_1B000000,
        64'h1E000000_03000000,
        64'h01000000_83000000,
        64'h04000000_03000000,
        64'h00000000_00000000,
        64'h04000000_03000000,
        64'h00000000_30303030,
        64'h30306340_72656C6C,
        64'h6F72746E_6F632D74,
        64'h70757272_65746E69,
        64'h01000000_02000000,
        64'h006C6F72_746E6F63,
        64'hD2000000_08000000,
        64'h03000000_00000C00,
        64'h00000000_00000002,
        64'h00000000_5B000000,
        64'h10000000_03000000,
        64'h07000000_01000000,
        64'h03000000_01000000,
        64'hBE000000_10000000,
        64'h03000000_00000000,
        64'h30746E69_6C632C76,
        64'h63736972_1B000000,
        64'h0D000000_03000000,
        64'h00000030_30303030,
        64'h30324074_6E696C63,
        64'h01000000_B7000000,
        64'h00000000_03000000,
        64'h00007375_622D656C,
        64'h706D6973_00636F73,
        64'h2D657261_622D656E,
        64'h61697261_2C687465,
        64'h1B000000_1F000000,
        64'h03000000_02000000,
        64'h0F000000_04000000,
        64'h03000000_02000000,
        64'h00000000_04000000,
        64'h03000000_00636F73,
        64'h01000000_02000000,
        64'h00000008_00000000,
        64'h00000080_00000000,
        64'h5B000000_10000000,
        64'h03000000_00007972,
        64'h6F6D656D_4F000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6F6D656D,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h01000000_AF000000,
        64'h04000000_03000000,
        64'h01000000_A9000000,
        64'h04000000_03000000,
        64'h00006374_6E692D75,
        64'h70632C76_63736972,
        64'h1B000000_0F000000,
        64'h03000000_94000000,
        64'h00000000_03000000,
        64'h01000000_83000000,
        64'h04000000_03000000,
        64'h00000000_72656C6C,
        64'h6F72746E_6F632D74,
        64'h70757272_65746E69,
        64'h01000000_79000000,
        64'h00000000_03000000,
        64'h40787D01_2C000000,
        64'h04000000_03000000,
        64'h00003933_76732C76,
        64'h63736972_70000000,
        64'h0B000000_03000000,
        64'h00007573_63616D69,
        64'h34367672_66000000,
        64'h0B000000_03000000,
        64'h00000076_63736972,
        64'h00656E61_69726120,
        64'h2C687465_1B000000,
        64'h12000000_03000000,
        64'h00000000_79616B6F,
        64'h5F000000_05000000,
        64'h03000000_00000000,
        64'h5B000000_04000000,
        64'h03000000_00757063,
        64'h4F000000_04000000,
        64'h03000000_00000000,
        64'h3F000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787D01_2C000000,
        64'h04000000_03000000,
        64'h00000000_0F000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_00657261,
        64'h622D656E_61697261,
        64'h2C687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2D657261,
        64'h622D656E_61697261,
        64'h2C687465_1B000000,
        64'h14000000_03000000,
        64'h02000000_0F000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h5C050000_47010000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h94050000_38000000,
        64'hDB060000_EDFE0DD0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_0000BFF5,
        64'h10500073_03C58593,
        64'h00000597_F1402573,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00008402_07458593,
        64'h00000597_F1402573,
        64'h01F41413_0010041B
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
