/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 835;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h0a0d2165_6e6f6420,
        64'h00000000_00206567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f63,
        64'h00000000_00000009,
        64'h3a656d61_6e090a0d,
        64'h00093a73_65747562,
        64'h69727474_61090a0d,
        64'h00000009_3a61626c,
        64'h20747361_6c090a0d,
        64'h0000093a_61626c20,
        64'h74737269_66090a0d,
        64'h00000000_00000000,
        64'h09202020_20203a64,
        64'h69756720_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_00000000,
        64'h093a6469_75672065,
        64'h70797420_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20747067,
        64'h00000009_20203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20657a69_73090a0d,
        64'h00000009_3a736569,
        64'h72746e65_206e6f69,
        64'h74697472_61702072,
        64'h65626d75_6e090a0d,
        64'h00000009_2020203a,
        64'h61626c20_73656972,
        64'h746e6520_6e6f6974,
        64'h69747261_70090a0d,
        64'h00093a61_646c2070,
        64'h756b6361_62090a0d,
        64'h00000000_00000000,
        64'h093a6162_6c20746e,
        64'h65727275_63090a0d,
        64'h00000009_3a646576,
        64'h72657365_72090a0d,
        64'h00093a72_65646165,
        64'h685f6372_63090a0d,
        64'h00000000_00000909,
        64'h3a657a69_73090a0d,
        64'h00000009_3a6e6f69,
        64'h73697665_72090a0d,
        64'h0000093a_65727574,
        64'h616e6769_73090a0d,
        64'h00000000_003a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20747067,
        64'h0000203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_63206473,
        64'h00000000_0000000a,
        64'h0d216465_7a696c61,
        64'h6974696e_69206473,
        64'h00000000_0a0d676e,
        64'h69746978_65202e2e,
        64'h2e647320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f63,
        64'h00000000_0000002e,
        64'h0000000a_0d202e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e69,
        64'h00000031_34646d63,
        64'h00000035_35646d63,
        64'h00000000_30646d63,
        64'h00000020_3a206573,
        64'h6e6f7073_65720920,
        64'h00000000_0020646e,
        64'h616d6d6f_63204453,
        64'h00000000_00000a0d,
        64'h65736e6f_70736572,
        64'h20647320_64696c61,
        64'h7620646e_69662074,
        64'h6f6e2064_6c756f63,
        64'h00000000_203f3f79,
        64'h74706d65_20746f6e,
        64'h206f6669_66207872,
        64'h00000000_00000a0d,
        64'h2164657a_696c6169,
        64'h74696e69_20495053,
        64'h00000000_00007830,
        64'h203a7375_74617473,
        64'h00000000_00000a0d,
        64'h49505320_74696e69,
        64'h00000a0d_21646c72,
        64'h6f57206f_6c6c6548,
        64'h00000000_0000006f,
        64'h69646d2d_7361682c,
        64'h786e6c78_006c616e,
        64'h7265746e_692d6573,
        64'h752c786e_6c780067,
        64'h6e6f702d_676e6970,
        64'h2d78742c_786e6c78,
        64'h00687464_69772d64,
        64'h692d6978_612d732c,
        64'h786e6c78_00676e6f,
        64'h702d676e_69702d78,
        64'h722c786e_6c780065,
        64'h636e6174_736e692c,
        64'h786e6c78_006f6964,
        64'h6d2d6564_756c636e,
        64'h692c786e_6c78006b,
        64'h63616270_6f6f6c2d,
        64'h6c616e72_65746e69,
        64'h2d656475_6c636e69,
        64'h2c786e6c_78007372,
        64'h65666675_622d6c61,
        64'h626f6c67_2d656475,
        64'h6c636e69_2c786e6c,
        64'h78007865_6c707564,
        64'h2c786e6c_7800656c,
        64'h646e6168_2d796870,
        64'h00737365_72646461,
        64'h2d63616d_2d6c6163,
        64'h6f6c0070_772d656c,
        64'h62617369_64007365,
        64'h676e6172_2d656761,
        64'h746c6f76_0079636e,
        64'h65757165_72662d78,
        64'h616d2d69_7073006f,
        64'h69746172_2d6b6373,
        64'h2c786e6c_78007374,
        64'h69622d72_6566736e,
        64'h6172742d_6d756e2c,
        64'h786e6c78_00737469,
        64'h622d7373_2d6d756e,
        64'h2c786e6c_78007473,
        64'h6978652d_6f666966,
        64'h2c786e6c_7800796c,
        64'h696d6166_2c786e6c,
        64'h78006874_6469772d,
        64'h6f692d67_65720074,
        64'h66696873_2d676572,
        64'h00737470_75727265,
        64'h746e6900_746e6572,
        64'h61702d74_70757272,
        64'h65746e69_00646565,
        64'h70732d74_6e657272,
        64'h75630076_65646e2c,
        64'h76637369_72007974,
        64'h69726f69_72702d78,
        64'h616d2c76_63736972,
        64'h0073656d_616e2d67,
        64'h65720064_65646e65,
        64'h7478652d_73747075,
        64'h72726574_6e690073,
        64'h65676e61_7200656c,
        64'h646e6168_702c7875,
        64'h6e696c00_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h02000000_02000000,
        64'h03000000_bb000000,
        64'h04000000_03000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h01000000_67000000,
        64'h04000000_03000000,
        64'h00000000_7968702d,
        64'h74656e72_65687465,
        64'h5b000000_0d000000,
        64'h03000000_00000000,
        64'h35313963_2e633130,
        64'h3064692d_7968702d,
        64'h74656e72_65687465,
        64'h1b000000_19000000,
        64'h03000000_00003040,
        64'h7968702d_74656e72,
        64'h65687465_01000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_6f69646d,
        64'h01000000_01000000,
        64'h94020000_04000000,
        64'h03000000_00000000,
        64'h82020000_04000000,
        64'h03000000_01000000,
        64'h70020000_04000000,
        64'h03000000_04000000,
        64'h5c020000_04000000,
        64'h03000000_01000000,
        64'h4a020000_04000000,
        64'h03000000_00657469,
        64'h6c74656e_72656874,
        64'h655f6978_615f786e,
        64'h6c785f69_3c020000,
        64'h18000000_03000000,
        64'h01000000_2a020000,
        64'h04000000_03000000,
        64'h00000000_0b020000,
        64'h04000000_03000000,
        64'h01000000_ef010000,
        64'h04000000_03000000,
        64'h01000000_e3010000,
        64'h04000000_03000000,
        64'h00000100_00000000,
        64'h00000030_00000000,
        64'h67000000_10000000,
        64'h03000000_03000000,
        64'hd8010000_04000000,
        64'h03000000_00002201,
        64'h00350a00_c6010000,
        64'h06000000_03000000,
        64'h00000000_03000000,
        64'h25010000_08000000,
        64'h03000000_02000000,
        64'h14010000_04000000,
        64'h03000000_006b726f,
        64'h7774656e_5b000000,
        64'h08000000_03000000,
        64'h0000612e_30302e31,
        64'h2d657469_6c74656e,
        64'h72656874_652d7370,
        64'h782c786e_6c780030,
        64'h2e332d65_74696c74,
        64'h656e7265_6874652d,
        64'h6978612c_786e6c78,
        64'h1b000000_37000000,
        64'h03000000_00000030,
        64'h30303030_30303340,
        64'h74656e72_65687465,
        64'h01000000_02000000,
        64'h02000000_bb010000,
        64'h00000000_03000000,
        64'he40c0000_e40c0000,
        64'hac010000_08000000,
        64'h03000000_20bcbe00,
        64'h9a010000_04000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00000000,
        64'h746f6c73_2d697073,
        64'h2d636d6d_1b000000,
        64'h0d000000_03000000,
        64'h00000030_40636d6d,
        64'h01000000_04000000,
        64'h8b010000_04000000,
        64'h03000000_08000000,
        64'h74010000_04000000,
        64'h03000000_01000000,
        64'h63010000_04000000,
        64'h03000000_01000000,
        64'h53010000_04000000,
        64'h03000000_00377865,
        64'h746e696b_47010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000020_00000000,
        64'h67000000_10000000,
        64'h03000000_02000000,
        64'h02000000_25010000,
        64'h08000000_03000000,
        64'h02000000_14010000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00612e30_302e322d,
        64'h6970732d_7370782c,
        64'h786e6c78_00622e30,
        64'h302e322d_6970732d,
        64'h7370782c_786e6c78,
        64'h1b000000_28000000,
        64'h03000000_00000000,
        64'h30303030_30303032,
        64'h40697073_2d737078,
        64'h01000000_02000000,
        64'h04000000_3a010000,
        64'h04000000_03000000,
        64'h02000000_30010000,
        64'h04000000_03000000,
        64'h01000000_25010000,
        64'h04000000_03000000,
        64'h02000000_14010000,
        64'h04000000_03000000,
        64'h00c20100_06010000,
        64'h04000000_03000000,
        64'h80f0fa02_4b000000,
        64'h04000000_03000000,
        64'h00100000_00000000,
        64'h00000010_00000000,
        64'h67000000_10000000,
        64'h03000000_00303537,
        64'h3631736e_1b000000,
        64'h08000000_03000000,
        64'h00000030_30303030,
        64'h30303140_74726175,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'hde000000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000000,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'hffff0000_01000000,
        64'hca000000_08000000,
        64'h03000000_00333130,
        64'h2d677562_65642c76,
        64'h63736972_1b000000,
        64'h10000000_03000000,
        64'h00003040_72656c6c,
        64'h6f72746e_6f632d67,
        64'h75626564_01000000,
        64'h02000000_02000000,
        64'hbb000000_04000000,
        64'h03000000_02000000,
        64'hb5000000_04000000,
        64'h03000000_03000000,
        64'hfb000000_04000000,
        64'h03000000_07000000,
        64'he8000000_04000000,
        64'h03000000_00000004,
        64'h00000000_0000000c,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h09000000_01000000,
        64'h0b000000_01000000,
        64'hca000000_10000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h00306369_6c702c76,
        64'h63736972_1b000000,
        64'h0c000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_00000000,
        64'h04000000_03000000,
        64'h00000000_30303030,
        64'h30306340_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'hde000000_08000000,
        64'h03000000_00000c00,
        64'h00000000_00000002,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h07000000_01000000,
        64'h03000000_01000000,
        64'hca000000_10000000,
        64'h03000000_00000000,
        64'h30746e69_6c632c76,
        64'h63736972_1b000000,
        64'h0d000000_03000000,
        64'h00000030_30303030,
        64'h30324074_6e696c63,
        64'h01000000_c3000000,
        64'h00000000_03000000,
        64'h00007375_622d656c,
        64'h706d6973_00636f73,
        64'h2d657261_622d656e,
        64'h61697261_2c687465,
        64'h1b000000_1f000000,
        64'h03000000_02000000,
        64'h0f000000_04000000,
        64'h03000000_02000000,
        64'h00000000_04000000,
        64'h03000000_00636f73,
        64'h01000000_02000000,
        64'h00000008_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h01000000_bb000000,
        64'h04000000_03000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00007573_63616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hf8080000_a2020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h30090000_38000000,
        64'hd20b0000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_a0018402,
        64'h02058593_00000597,
        64'h01f41413_0010041b,
        64'hd71ff0ef_057e65a1,
        64'h4505f58f_f0efc165,
        64'h05130000_1517f32f,
        64'hf0efe406_1141bb75,
        64'h8156f70f_f0eff0e5,
        64'h05130000_1517c75f,
        64'hf0ef855a_865e020a,
        64'h2583f88f_f0eff0e5,
        64'h05130000_1517f589,
        64'h93e30804_8493f9cf,
        64'hf0ef2985_c9c50513,
        64'h00001517_ff2c9be3,
        64'h873ff0ef_09050009,
        64'h4503fb8f_f0eff2e5,
        64'h05130000_1517847f,
        64'hf0ef7088_fcaff0ef,
        64'hf3050513_00001517,
        64'h859ff0ef_6c88fdcf,
        64'hf0eff325_05130000,
        64'h151786bf_f0ef0704,
        64'h8c930284_89136888,
        64'hff6ff0ef_f3c50513,
        64'h00001517_ff991be3,
        64'h8cbff0ef_09050009,
        64'h45030109_0c93815f,
        64'hf0eff3a5_05130000,
        64'h1517fe99_1be38e9f,
        64'hf0ef0905_00094503,
        64'hff048913_833ff0ef,
        64'hf3850513_00001517,
        64'h903ff0ef_0ff9f513,
        64'h847ff0ef_f3450513,
        64'h00001517_4c11010a,
        64'h0493859f_f0efd565,
        64'h05130000_15178e7f,
        64'hf0ef8526_86bff0ef,
        64'he4850513_00001517,
        64'hc10584aa_8a0ad75f,
        64'hf0ef850a_46057101,
        64'h44ac889f_f0efd865,
        64'h05130000_15178d7f,
        64'hf0ef48e8_89bff0ef,
        64'hf6850513_00001517,
        64'h8e9ff0ef_48a88adf,
        64'hf0eff5a5_05130000,
        64'h151793bf_f0ef64a8,
        64'h8bfff0ef_f4c50513,
        64'h00001517_94dff0ef,
        64'h70888d1f_f0eff4e5,
        64'h05130000_151795ff,
        64'hf0ef6c88_8e3ff0ef,
        64'hf4850513_00001517,
        64'h931ff0ef_48c88f5f,
        64'hf0eff4a5_05130000,
        64'h1517943f_f0ef4888,
        64'h907ff0ef_f4c50513,
        64'h00001517_955ff0ef,
        64'h44c8919f_f0eff4e5,
        64'h05130000_1517967f,
        64'hf0ef4488_92bff0ef,
        64'hf5050513_00001517,
        64'h9b9ff0ef_608893df,
        64'hf0eff525_05130000,
        64'h1517949f_f0eff3e5,
        64'h05130000_1517955f,
        64'hf0efe525_05130000,
        64'h15179e3f_f0ef854a,
        64'h967ff0ef_f4450513,
        64'h00001517_c105892a,
        64'h848ae71f_f0ef850a,
        64'h45854605_71018a8a,
        64'h987ff0ef_f4c50513,
        64'h00001517_89aa8082,
        64'h61256ca2_6c426be2,
        64'h7b027aa2_7a4279e2,
        64'h690664a6_644660e6,
        64'hfa040113_9b3ff0ef,
        64'hf5050513_00001517,
        64'hc515e1df_f0ef8bae,
        64'h8b2a1080_e466e862,
        64'hf456f852_fc4ee0ca,
        64'he4a6ec86_ec5ef05a,
        64'he8a2711d_bfe15479,
        64'h80826169_6baa6b4a,
        64'h6aea7a0a_79aa794a,
        64'h74ea640e_60ae8522,
        64'hc79ff0ef_c85ff0ef,
        64'h45314581_46054401,
        64'hf89046e3_14fda15f,
        64'hf0effaa5_05130000,
        64'h1517e799_0354e7b3,
        64'h05341263_29819041,
        64'h14428c49_cadff0ef,
        64'h90410305_14138922,
        64'h0085151b_cbdff0ef,
        64'hfd641ae3_04040413,
        64'hff7917e3_89aaf0ff,
        64'hf0ef0905_854e0007,
        64'hc5830124_07b30400,
        64'h0b934901_c65ff0ef,
        64'h850a0400_05938622,
        64'h4981844a_20090b13,
        64'hff451ee3_cfdff0ef,
        64'h3e800a93_0fe00a13,
        64'h90811482_bff5d0ff,
        64'hf0efc501_d1dff0ef,
        64'h454985a2_0ff67613,
        64'h00166613_0015161b,
        64'hf4fff0ef_0ff47593,
        64'hf57ff0ef_0ff5f593,
        64'h0084559b_f63ff0ef,
        64'h0ff5f593_0104559b,
        64'hf6fff0ef_45010ff5,
        64'hf5930184_559bfee7,
        64'h9be30785_00c68023,
        64'h00f106b3_08000713,
        64'h567d4781_842e892a,
        64'he55ee95a_ed56f152,
        64'hf54ee586_84b2f94a,
        64'hfd26e1a2_71558082,
        64'h91411542_8d3d8ff9,
        64'h0057979b_17016709,
        64'h0107d79b_0105179b,
        64'h4105551b_0105151b,
        64'h8d2d00c5_95138da9,
        64'h893d0045_d51b8da9,
        64'h91411542_8d5d0522,
        64'h0085579b_808207f5,
        64'h75138d2d_00451593,
        64'h8d2d8d3d_0045d51b,
        64'h0075d79b_8de98082,
        64'h0141853e_640260a2,
        64'h4781c111_57f5f89f,
        64'hf0efc511_57f9efbf,
        64'hf0efc911_57fdec9f,
        64'hf0effc6d_e05ff0ef,
        64'h347d4429_b93ff0ef,
        64'h11050513_00001517,
        64'hc8bff0ef_e022e406,
        64'h11418082_61050015,
        64'h351364a2_644260e2,
        64'h0004051b_fc940ce3,
        64'he39ff0ef_ec5ff0ef,
        64'h13850513_00001517,
        64'h85aa842a_e55ff0ef,
        64'h02900513_400005b7,
        64'h07700613_fbdff0ef,
        64'h4485e822_ec06e426,
        64'h11018082_01410015,
        64'h3513157d_640260a2,
        64'h0004051b_f05ff0ef,
        64'h17250513_85a20000,
        64'h1517e8bf_f0ef842a,
        64'he99ff0ef_e022e406,
        64'h03700513_45810650,
        64'h06131141_80826105,
        64'h690264a2_644260e2,
        64'h00153513_f5650513,
        64'h0004051b_01249863,
        64'h88bd00f9_1b634501,
        64'h4785ecbf_f0efecff,
        64'hf0ef842a_ed5ff0ef,
        64'h84aaedbf_f0efedff,
        64'hf0efee3f_f0ef892a,
        64'hef1ff0ef_e04ae426,
        64'he822ec06_45211aa0,
        64'h05930870_06131101,
        64'h80826105_450564a2,
        64'h644260e2_fe9410e3,
        64'hf99ff0ef_1fe50513,
        64'h85a20000_1517f1ff,
        64'hf0ef842a_f2dff0ef,
        64'h45010950_06134581,
        64'h4485e822_ec06e426,
        64'h1101cc1f_f06f6105,
        64'h1c050513_00001517,
        64'h60e26442_d97ff0ef,
        64'h852e65a2_cdbff0ef,
        64'h23050513_00001517,
        64'hce7ff0ef_8522cedf,
        64'hf0efe42e_ec062365,
        64'h05130000_1517842a,
        64'he8221101_80826145,
        64'h64e28526_740270a2,
        64'hd0fff0ef_22c50513,
        64'h00001517_f475147d,
        64'h0007da63_84aa4187,
        64'hd79b0185_179bfa7f,
        64'hf0efeb5f_f0ef8532,
        64'h06400413_6622ec1f,
        64'hf0ef0ff4_7513ec9f,
        64'hf0ef0ff5_75130084,
        64'h551bed5f_f0ef0ff5,
        64'h75130104_551bee1f,
        64'hf0ef0ff5_75130184,
        64'h551beedf_f0ef0404,
        64'he513febf_f0ef84aa,
        64'h842eec26_f022e432,
        64'hf4067179_f07ff06f,
        64'h0ff00513_8082557d,
        64'hb7e900d7_00230785,
        64'h00f60733_06c82683,
        64'hff798b05_5178bf4d,
        64'hd6b80785_0007c703,
        64'h80824501_d3b84719,
        64'hdbb8577d_200007b7,
        64'h00b6ef63_0007869b,
        64'h20000837_20000537,
        64'hfff58b85_537c2000,
        64'h0737d3b8_200007b7,
        64'h10600713_fff537fd,
        64'h00010320_079304b7,
        64'h616340a7_873b87aa,
        64'h200006b7_dbb85779,
        64'h200007b7_06b7ec63,
        64'h10000793_80826105,
        64'h64a2d3b8_4719dbb8,
        64'h644260e2_0ff47513,
        64'h577d2000_07b7e25f,
        64'hf0ef3225_05130000,
        64'h1517eb3f_f0ef9101,
        64'h15024088_e3bff0ef,
        64'h34050513_00001517,
        64'he3958b85_240153fc,
        64'h57e0ff65_8b050647,
        64'h849353f8_d3b81060,
        64'h07132000_07b7fff5,
        64'h37fd0001_06400793,
        64'hd7a8dbb8_5779e426,
        64'he822ec06_200007b7,
        64'h1101e81f_f06f6105,
        64'h37050513_00001517,
        64'h64a260e2_6442d03c,
        64'h4799e99f_f0ef3965,
        64'h05130000_1517f27f,
        64'hf0ef9101_02049513,
        64'h2481eb1f_f0ef38e5,
        64'h05130000_15175064,
        64'hd03c1660_0793ec5f,
        64'hf0ef3c25_05130000,
        64'h1517f53f_f0ef9101,
        64'h02049513_2481eddf,
        64'hf0ef3ba5_05130000,
        64'h15175064_d03c1040,
        64'h07932000_0437fff5,
        64'h37fd0001_47a9c3b8,
        64'h47292000_07b7f05f,
        64'hf0efe426_e822ec06,
        64'h3da50513_11010000,
        64'h15178082_41088082,
        64'hc10c8082_610560e2,
        64'hee1ff0ef_00914503,
        64'hee9ff0ef_00814503,
        64'hf55ff0ef_ec06002c,
        64'h11018082_61456942,
        64'h64e27402_70a2fe94,
        64'h10e3f0bf_f0ef0091,
        64'h4503f13f_f0ef3461,
        64'h00814503_f81ff0ef,
        64'h0ff57513_002c0089,
        64'h553354e1_03800413,
        64'h892af406_e84aec26,
        64'hf0227179_80826145,
        64'h694264e2_740270a2,
        64'hfe9410e3_f4dff0ef,
        64'h00914503_f55ff0ef,
        64'h34610081_4503fc3f,
        64'hf0ef0ff5_7513002c,
        64'h0089553b_54e14461,
        64'h892af406_e84aec26,
        64'hf0227179_808200f5,
        64'h80230007_c78300e5,
        64'h80a397aa_81110007,
        64'h4703973e_00f57713,
        64'h88078793_00002797,
        64'hb7f50405_fa5ff0ef,
        64'h80820141_640260a2,
        64'he5090004_4503842a,
        64'he406e022_11418082,
        64'h00e78823_02000713,
        64'h00e78423_fc700713,
        64'h00e78623_470d0007,
        64'h822300e7_8023476d,
        64'h00e78623_f8000713,
        64'h00078223_100007b7,
        64'h808200a7_0023dfe5,
        64'h0207f793_01474783,
        64'h10000737_80820205,
        64'h75130147_c5031000,
        64'h07b78082_00054503,
        64'h808200b5_00238082,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_01f49493,
        64'h0010049b_9c458593,
        64'h00001597_f1402573,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'hfe091ee3_0004a903,
        64'h00092023_00990933,
        64'h00291913_f1402973,
        64'h020004b7_fe090ae3,
        64'h00897913_34402973,
        64'h10500073_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_0124a023,
        64'h00100913_020004b7,
        64'h1df000ef_01a11113,
        64'h0210011b_03249663,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
