`define ARTY_A7_100

`define ARIANE_DATA_WIDTH 64

// Instantiate protocl checker
// `define PROTOCOL_CHECKER

// write-back cache
// `define WB_DCACHE

// write-through cache
`define WT_DCACHE

// causes build error in cdc_2phase_clearable.sv
`define COMMON_CELLS_ASSERTS_OFF

`define RAMB16
