/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 911;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'h0a0d2165_6e6f6420,
        64'h00000000_00206567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f63,
        64'h00000000_00000009,
        64'h3a656d61_6e090a0d,
        64'h00093a73_65747562,
        64'h69727474_61090a0d,
        64'h00000009_3a61626c,
        64'h20747361_6c090a0d,
        64'h0000093a_61626c20,
        64'h74737269_66090a0d,
        64'h00000000_00000000,
        64'h09202020_20203a64,
        64'h69756720_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_00000000,
        64'h093a6469_75672065,
        64'h70797420_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20747067,
        64'h00000009_20203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20657a69_73090a0d,
        64'h00000009_3a736569,
        64'h72746e65_206e6f69,
        64'h74697472_61702072,
        64'h65626d75_6e090a0d,
        64'h00000009_2020203a,
        64'h61626c20_73656972,
        64'h746e6520_6e6f6974,
        64'h69747261_70090a0d,
        64'h00093a61_646c2070,
        64'h756b6361_62090a0d,
        64'h00000000_00000000,
        64'h093a6162_6c20746e,
        64'h65727275_63090a0d,
        64'h00000009_3a646576,
        64'h72657365_72090a0d,
        64'h00093a72_65646165,
        64'h685f6372_63090a0d,
        64'h00000000_00000909,
        64'h3a657a69_73090a0d,
        64'h00000009_3a6e6f69,
        64'h73697665_72090a0d,
        64'h0000093a_65727574,
        64'h616e6769_73090a0d,
        64'h00000000_003a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20747067,
        64'h0000203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_63206473,
        64'h00000000_0000000a,
        64'h0d216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_0000000a,
        64'h0d216465_7a696c61,
        64'h6974696e_69206473,
        64'h00000000_0a0d676e,
        64'h69746978_65202e2e,
        64'h2e647320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f63,
        64'h00000000_0000002e,
        64'h00000000_0000000a,
        64'h0d6b636f_6c622044,
        64'h53206461_65722074,
        64'h6f6e2064_6c756f63,
        64'h0000000a_0d202e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e69,
        64'h00000031_34646d63,
        64'h00000035_35646d63,
        64'h00000000_30646d63,
        64'h00000020_3a206573,
        64'h6e6f7073_65720920,
        64'h00000000_0020646e,
        64'h616d6d6f_63204453,
        64'h00000000_203f3f79,
        64'h74706d65_20746f6e,
        64'h206f6669_66207872,
        64'h00000000_00000a0d,
        64'h2164657a_696c6169,
        64'h74696e69_20495053,
        64'h00000000_00007830,
        64'h203a7375_74617473,
        64'h00000000_00000a0d,
        64'h49505320_74696e69,
        64'h00000000_0000000a,
        64'h0a0a0a0d_21646c72,
        64'h6f57206f_6c6c6548,
        64'h00000000_00000032,
        64'h2d746c75_61666564,
        64'h2d697274_2c786e6c,
        64'h7800746c_75616665,
        64'h642d6972_742c786e,
        64'h6c78006c_6175642d,
        64'h73692c78_6e6c7800,
        64'h746e6573_6572702d,
        64'h74707572_7265746e,
        64'h692c786e_6c780068,
        64'h74646977_2d326f69,
        64'h70672c78_6e6c7800,
        64'h68746469_772d6f69,
        64'h70672c78_6e6c7800,
        64'h322d746c_75616665,
        64'h642d7475_6f642c78,
        64'h6e6c7800_746c7561,
        64'h6665642d_74756f64,
        64'h2c786e6c_7800322d,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h72656c6c_6f72746e,
        64'h6f632d6f_69706700,
        64'h736c6c65_632d6f69,
        64'h70672300_73736572,
        64'h6464612d_63616d2d,
        64'h6c61636f_6c007077,
        64'h2d656c62_61736964,
        64'h00736567_6e61722d,
        64'h65676174_6c6f7600,
        64'h79636e65_75716572,
        64'h662d7861_6d2d6970,
        64'h73006f69_7461722d,
        64'h6b63732c_786e6c78,
        64'h00737469_622d7265,
        64'h66736e61_72742d6d,
        64'h756e2c78_6e6c7800,
        64'h73746962_2d73732d,
        64'h6d756e2c_786e6c78,
        64'h00747369_78652d6f,
        64'h6669662c_786e6c78,
        64'h00796c69_6d61662c,
        64'h786e6c78_00687464,
        64'h69772d6f_692d6765,
        64'h72007466_6968732d,
        64'h67657200_73747075,
        64'h72726574_6e690074,
        64'h6e657261_702d7470,
        64'h75727265_746e6900,
        64'h64656570_732d746e,
        64'h65727275_63007665,
        64'h646e2c76_63736972,
        64'h00797469_726f6972,
        64'h702d7861_6d2c7663,
        64'h73697200_73656d61,
        64'h6e2d6765_72006465,
        64'h646e6574_78652d73,
        64'h74707572_7265746e,
        64'h69007365_676e6172,
        64'h00646564_6e657073,
        64'h75732d65_74617473,
        64'h2d6e6961_74657200,
        64'h72656767_6972742d,
        64'h746c7561_6665642c,
        64'h78756e69_6c00736f,
        64'h69706700_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'hffffffff_bf020000,
        64'h04000000_03000000,
        64'hffffffff_ae020000,
        64'h04000000_03000000,
        64'h01000000_a1020000,
        64'h04000000_03000000,
        64'h00000000_8a020000,
        64'h04000000_03000000,
        64'h08000000_79020000,
        64'h04000000_03000000,
        64'h08000000_69020000,
        64'h04000000_03000000,
        64'h00000000_55020000,
        64'h04000000_03000000,
        64'h00000000_43020000,
        64'h04000000_03000000,
        64'h00000000_31020000,
        64'h04000000_03000000,
        64'h00000000_21020000,
        64'h04000000_03000000,
        64'h00000100_00000000,
        64'h00000040_00000000,
        64'h67000000_10000000,
        64'h03000000_11020000,
        64'h00000000_03000000,
        64'h00000000_612e3030,
        64'h2e312d6f_6970672d,
        64'h7370782c_786e6c78,
        64'h1b000000_15000000,
        64'h03000000_02000000,
        64'h05020000_04000000,
        64'h03000000_00000030,
        64'h30303030_30303440,
        64'h6f697067_01000000,
        64'h02000000_00800000,
        64'h00000000_00000030,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00007fe3_023e1800,
        64'hf3010000_06000000,
        64'h03000000_00000000,
        64'h03000000_52010000,
        64'h08000000_03000000,
        64'h03000000_41010000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_00687465,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_00000000,
        64'h30303030_30303033,
        64'h40687465_2d637369,
        64'h72776f6c_01000000,
        64'h02000000_02000000,
        64'he8010000_00000000,
        64'h03000000_e40c0000,
        64'he40c0000_d9010000,
        64'h08000000_03000000,
        64'h20bcbe00_c7010000,
        64'h04000000_03000000,
        64'h00000000_67000000,
        64'h04000000_03000000,
        64'h00000000_746f6c73,
        64'h2d697073_2d636d6d,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h40636d6d_01000000,
        64'h04000000_b8010000,
        64'h04000000_03000000,
        64'h08000000_a1010000,
        64'h04000000_03000000,
        64'h01000000_90010000,
        64'h04000000_03000000,
        64'h01000000_80010000,
        64'h04000000_03000000,
        64'h00377865_746e696b,
        64'h74010000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h02000000_02000000,
        64'h52010000_08000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_00612e30,
        64'h302e322d_6970732d,
        64'h7370782c_786e6c78,
        64'h00622e30_302e322d,
        64'h6970732d_7370782c,
        64'h786e6c78_1b000000,
        64'h28000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40697073,
        64'h2d737078_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h03000000_41010000,
        64'h04000000_03000000,
        64'h00100000_00000000,
        64'h00000018_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h06000000_05000000,
        64'h04000000_52010000,
        64'h10000000_03000000,
        64'h00007265_6d69745f,
        64'h6270612c_706c7570,
        64'h1b000000_0f000000,
        64'h03000000_00003030,
        64'h30303030_38314072,
        64'h656d6974_01000000,
        64'h02000000_04000000,
        64'h67010000_04000000,
        64'h03000000_02000000,
        64'h5d010000_04000000,
        64'h03000000_01000000,
        64'h52010000_04000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00c20100,
        64'h33010000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000010,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00303537_3631736e,
        64'h1b000000_08000000,
        64'h03000000_00000030,
        64'h30303030_30303140,
        64'h74726175_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000000_00000000,
        64'h67000000_10000000,
        64'h03000000_ffff0000,
        64'h02000000_f7000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00003040,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h1e000000_28010000,
        64'h04000000_03000000,
        64'h07000000_15010000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h02000000_0b000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hf0000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_02000000,
        64'hd9000000_00000000,
        64'h03000000_00000074,
        64'h61656274_72616568,
        64'hc3000000_0a000000,
        64'h03000000_00000000,
        64'h01000000_01000000,
        64'hbd000000_0c000000,
        64'h03000000_00000064,
        64'h656c2d74_61656274,
        64'h72616568_01000000,
        64'h00000073_64656c2d,
        64'h6f697067_1b000000,
        64'h0a000000_03000000,
        64'h00000000_7364656c,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'hc0e1e400_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h60090000_d2020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h98090000_38000000,
        64'h6a0c0000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_0000bf61,
        64'hdc6ff0ef_10000537,
        64'hfff44583_dd2ff0ef,
        64'h10000537_ffe44583,
        64'hddeff0ef_10000537,
        64'hffd44583_deaff0ef,
        64'h04111000_05370004,
        64'h4583a001_dfaff0ef,
        64'h02050513_45811000,
        64'h0537fe94_17e3e2af,
        64'hf0ef0ff5_7513ff25,
        64'h0de3842a_f72ff0ef,
        64'h44b5597d_e28ff0ef,
        64'h10000537_02941b63,
        64'he60ff0ef_01440493,
        64'he04aec06_e426eb64,
        64'h04130805_05132005,
        64'h85930000_141702fa,
        64'hf53765f1_e8221101,
        64'hb38deccf_f0ef1c65,
        64'h05130000_1517bbd9,
        64'hf2050513_00001517,
        64'hf64ff0ef_8526ee8f,
        64'hf0ef0225_05130000,
        64'h1517ef4f_f0ef0165,
        64'h05130000_1517bbfd,
        64'hf4850513_00001517,
        64'hf8cff0ef_8526f10f,
        64'hf0ef04a5_05130000,
        64'h1517f1cf_f0ef03e5,
        64'h05130000_1517c929,
        64'h84aac3bf_f0ef8556,
        64'h865a020b_a583f38f,
        64'hf0ef21a5_05130000,
        64'h1517f384_9de30809,
        64'h0913080a_0993f50f,
        64'hf0ef2485_f9c50513,
        64'h00001517_ff3a1be3,
        64'h827ff0ef_0a05000a,
        64'h4503f6cf_f0ef23e5,
        64'h05130000_1517ffaf,
        64'hf0ef0109_3503f80f,
        64'hf0ef2425_05130000,
        64'h151780ff_f0ef0089,
        64'h3503f94f_f0ef2465,
        64'h05130000_1517823f,
        64'hf0effb89_8a130009,
        64'h3503facf_f0ef24e5,
        64'h05130000_1517ff2a,
        64'h1be3881f_f0ef0a05,
        64'h000a4503_f9098a13,
        64'hfcaff0ef_24c50513,
        64'h00001517_ff9a19e3,
        64'h89fff0ef_0a050007,
        64'hc503014d_07b34a01,
        64'hfeaff0ef_f8098d13,
        64'h25050513_00001517,
        64'h8bfff0ef_0ff4f513,
        64'h803ff0ef_24c50513,
        64'h00001517_4c114cc1,
        64'h10051b63_02010913,
        64'h08010993_84aa8b8a,
        64'hd31ff0ef_850a4605,
        64'h71010489_2583831f,
        64'hf0ef07a5_05130000,
        64'h151787ff_f0ef4556,
        64'h843ff0ef_26c50513,
        64'h00001517_891ff0ef,
        64'h4546855f_f0ef25e5,
        64'h05130000_15178e3f,
        64'hf0ef6526_867ff0ef,
        64'h25050513_00001517,
        64'h8f5ff0ef_7502879f,
        64'hf0ef2525_05130000,
        64'h1517907f_f0ef6562,
        64'h88bff0ef_24c50513,
        64'h00001517_8d9ff0ef,
        64'h455289df_f0ef24e5,
        64'h05130000_15178ebf,
        64'hf0ef4542_8afff0ef,
        64'h25050513_00001517,
        64'h8fdff0ef_45328c1f,
        64'hf0ef2525_05130000,
        64'h151790ff_f0ef4522,
        64'h8d3ff0ef_25450513,
        64'h00001517_961ff0ef,
        64'h65028e5f_f0ef2565,
        64'h05130000_15178f1f,
        64'hf0ef2425_05130000,
        64'h1517bf51_54f9901f,
        64'hf0ef14a5_05130000,
        64'h151798ff_f0ef8526,
        64'h913ff0ef_24c50513,
        64'h00001517_91fff0ef,
        64'h24050513_00001517,
        64'hc90584aa_890ae3ff,
        64'hf0ef850a_45854605,
        64'h710193df_f0ef2465,
        64'h05130000_15178082,
        64'h61256d02_6ca26c42,
        64'h6be27b02_7aa27a42,
        64'h79e26906_64a66446,
        64'h852660e6_fa040113,
        64'h54fd96df_f0ef24e5,
        64'h05130000_1517c90d,
        64'hdf1ff0ef_8b2e8aaa,
        64'h1080e06a_e466e862,
        64'hec5ef852_fc4ee0ca,
        64'he4a6ec86_f05af456,
        64'he8a2711d_b7655479,
        64'h80826169_6baa6b4a,
        64'h6aea7a0a_79aa794a,
        64'h74ea640e_852260ae,
        64'h547d9bdf_f0ef2765,
        64'h05130000_1517c5ff,
        64'hf0efc63f_f0efc67f,
        64'hf0efc6bf_f0efc6ff,
        64'hf0efc73f_f0efc77f,
        64'hf0efc7bf_f0efa805,
        64'hc81ff0ef_c8bff0ef,
        64'h45314581_46054401,
        64'hf93045e3_20048493,
        64'h19fda05f_f0ef2de5,
        64'h05130000_1517e799,
        64'h0359e7b3_07241c63,
        64'h29019041_14428c49,
        64'hcb9ff0ef_90411442,
        64'h0085141b_cc5ff0ef,
        64'hfc9418e3_04040413,
        64'hff7b15e3_892af19f,
        64'hf0ef0ff5_f5930b05,
        64'h854a0007_c5830164,
        64'h07b30400_0b934b01,
        64'hc6dff0ef_850a0400,
        64'h05938622_4901ff45,
        64'h1ee3d03f_f0efe004,
        64'h84133e80_0a930fe0,
        64'h0a13e959_20048493,
        64'hd1fff0ef_454985a2,
        64'h0ff67613_00166613,
        64'h00151613_f51ff0ef,
        64'h0ff47593_f59ff0ef,
        64'h0ff5f593_0084559b,
        64'hf65ff0ef_0ff5f593,
        64'h0104559b_f71ff0ef,
        64'h45010184_559bfee7,
        64'h9be30785_00c68023,
        64'h00f106b3_08000713,
        64'h567d4781_0209d993,
        64'h842e84aa_e55ee95a,
        64'hed56f152_f94ae586,
        64'hfd26e1a2_02061993,
        64'hf54e7155_80829141,
        64'h15428d2d_8d7d0055,
        64'h151b1781_67890105,
        64'h551b0105_951b8da9,
        64'h00c59513_8da9893d,
        64'h0045d51b_8da99141,
        64'h15428d5d_05220085,
        64'h579b8082_07f57513,
        64'h8d2d0045_15938d2d,
        64'h0ff57513_8d3d0045,
        64'hd51b0075_d79b8de9,
        64'h80820141_853e6402,
        64'h60a257f5_e1114781,
        64'hf89ff0ef_c51157f9,
        64'hefbff0ef_c91157fd,
        64'heb7ff0ef_fc6de07f,
        64'hf0ef347d_4429b79f,
        64'hf0ef41a5_05130000,
        64'h1517c8bf_f0efe022,
        64'he4061141_80826105,
        64'h00153513_64a26442,
        64'h0004051b_60e2fc94,
        64'h0ce3e3bf_f0efeb3f,
        64'hf0ef4425_05130000,
        64'h151785aa_842ae55f,
        64'hf0ef0290_05134000,
        64'h05b70770_0613fbdf,
        64'hf0ef4485_e822ec06,
        64'he4261101_80820141,
        64'h00153513_157d6402,
        64'h0004051b_60a2ef3f,
        64'hf0ef47c5_051385a2,
        64'h00001517_e8dff0ef,
        64'h842ae99f_f0efe022,
        64'he4060370_05134581,
        64'h06500613_11418082,
        64'h61056902_64a26442,
        64'h60e20015_3513f565,
        64'h05130004_051b0124,
        64'h986388bd_00f91b63,
        64'h45014785_ecdff0ef,
        64'hed1ff0ef_842aed7f,
        64'hf0ef84aa_eddff0ef,
        64'hee1ff0ef_ee5ff0ef,
        64'h892aef1f_f0efe04a,
        64'he426e822_ec064521,
        64'h1aa00593_08700613,
        64'h1101bfcd_45018082,
        64'h61056902_64a26442,
        64'h60e24505_f89ff0ef,
        64'h458550a5_05130000,
        64'h1517ff24_95e3c00d,
        64'hf29ff0ef_84aa347d,
        64'hf37ff0ef_45014581,
        64'h09500613_49057104,
        64'h0413e426_ec06e04a,
        64'h6409e822_1101b95d,
        64'h61055025_05130000,
        64'h151764a2_60e26442,
        64'hd8fff0ef_8522cd1f,
        64'hf0ef54a5_05130000,
        64'h1517cddf_f0ef8526,
        64'hce3ff0ef_842ee822,
        64'hec065525_05130000,
        64'h151784aa_e4261101,
        64'h80826105_690264a2,
        64'h644260e2_f47d147d,
        64'h0007d463_4187d79b,
        64'h0185179b_fadff0ef,
        64'h06400413_ebbff0ef,
        64'h8526ec1f_f0ef0ff4,
        64'h7513ec9f_f0ef0ff5,
        64'h75130084_551bed5f,
        64'hf0ef0ff5_75130104,
        64'h551bee1f_f0ef0184,
        64'h551bee9f_f0ef0409,
        64'h6513febf_f0ef892a,
        64'he04a84b2_842ee426,
        64'he822ec06_1101b709,
        64'h0ff00513_8082557d,
        64'hb7d900d7_00230785,
        64'h00f60733_06c82683,
        64'hff698b05_5178b77d,
        64'hd6b80785_00074703,
        64'h00f50733_80824501,
        64'hd3b84719_dbb8577d,
        64'h200007b7_02b6e163,
        64'h0007869b_20000837,
        64'h20000537_fff58b85,
        64'h537c2000_0737d3b8,
        64'h200007b7_10600713,
        64'hfff537fd_00010320,
        64'h079304b7_61630007,
        64'h871b4781_200006b7,
        64'hdbb85779_200007b7,
        64'h06b7ee63_10000793,
        64'h80826105_64a2d3b8,
        64'h4719dbb8_64420ff4,
        64'h7513577d_200007b7,
        64'h60e2e0df_f0ef6565,
        64'h05130000_1517e9bf,
        64'hf0ef9101_15024088,
        64'he23ff0ef_67450513,
        64'h00001517_e3958b85,
        64'h240153fc_57e0ff65,
        64'h8b050647_849353f8,
        64'hd3b81060_07132000,
        64'h07b7fff5_37fd0001,
        64'h06400793_d7a8dbb8,
        64'h5779e426_e822ec06,
        64'h200007b7_1101b59d,
        64'h61056a25_05130000,
        64'h151764a2_60e26442,
        64'hd03c4799_e7fff0ef,
        64'h6c850513_00001517,
        64'hf0dff0ef_91010204,
        64'h95132481_e97ff0ef,
        64'h6c050513_00001517,
        64'h5064d03c_16600793,
        64'heabff0ef_6f450513,
        64'h00001517_f39ff0ef,
        64'h91010204_95132481,
        64'hec3ff0ef_6ec50513,
        64'h00001517_5064d03c,
        64'h10400793_20000437,
        64'hfff537fd_000147a9,
        64'hc3b84729_200007b7,
        64'heebff0ef_e426e822,
        64'hec0670c5_05131101,
        64'h00001517_80822501,
        64'h41088082_c10c8082,
        64'h0ff57513_00074503,
        64'hc7898b85_557d0147,
        64'h47831000_07378082,
        64'h610560e2_ed1ff0ef,
        64'h00914503_ed9ff0ef,
        64'h00814503_f55ff0ef,
        64'hec06002c_11018082,
        64'h61456942_64e27402,
        64'h70a2ff24_10e3efbf,
        64'hf0ef0091_4503f03f,
        64'hf0ef3461_00814503,
        64'hf81ff0ef_0ff57513,
        64'h002c0084_d5335961,
        64'h03800413_84aaf406,
        64'he84aec26_f0227179,
        64'h80826145_694264e2,
        64'h740270a2_ff2410e3,
        64'hf3dff0ef_00914503,
        64'hf45ff0ef_34610081,
        64'h4503fc3f_f0ef0ff5,
        64'h7513002c_0084d53b,
        64'h59614461_84aaf406,
        64'he84aec26_f0227179,
        64'h808200f5_80230007,
        64'hc78300e5_80a397aa,
        64'h81110007_4703973e,
        64'h00f57713_a6c78793,
        64'h00001797_b7f50405,
        64'hf95ff0ef_80820141,
        64'h640260a2_e5090004,
        64'h4503842a_e406e022,
        64'h11418082_00e78823,
        64'h02000713_00e78423,
        64'h571d00e7_8623470d,
        64'h00a78223_0ff57513,
        64'h00e78023_0085551b,
        64'h0ff57713_00e78623,
        64'hf8000713_00078223,
        64'h100007b7_02b5553b,
        64'h0045959b_808200a7,
        64'h0023dfe5_0207f793,
        64'h01474783_10000737,
        64'h80820205_75130147,
        64'hc5031000_07b78082,
        64'h0ff57513_00054503,
        64'h808200b5_00238082,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_01f49493,
        64'h0010049b_c8458593,
        64'h00001597_f1402573,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'hfe091ee3_0004a903,
        64'h00092023_00990933,
        64'h00291913_f1402973,
        64'h020004b7_fe090ae3,
        64'h00897913_34402973,
        64'h10500073_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_0124a023,
        64'h00100913_020004b7,
        64'h295000ef_01a11113,
        64'h0210011b_03249663,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
